----------------------------------
--		Library Declaration 	--
----------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

----------------------------------
--		Entity Declaration 		--
----------------------------------

entity qft_2qbit is
	port(
		clk : in std_logic;
		reset : in std_logic; -- (Key0) on keypress, reset becomes zero, state becomes idle and input is taken. Press before start.
		start : in std_logic; -- (key1) on keypress, start becomes 0 and computation starts.
--		a0RE : in sfixed(4 downto -4); 
--		a1RE : in sfixed(4 downto -4);
--		a2RE : in sfixed(4 downto -4);
--		a3RE : in sfixed(4 downto -4);
--		a0IM : in sfixed(4 downto -4); 
--		a1IM : in sfixed(4 downto -4); 
--		a2IM : in sfixed(4 downto -4);
--		a3IM : in sfixed(4 downto -4);
--		b0RE : out sfixed(4 downto -4); -- first bit represents sign with remaining in 2s complement for negative number.
--		b1RE : out sfixed(4 downto -4); -- Actually only 8 out of 9 bits for storing data.
--		b2RE : out sfixed(4 downto -4);
--		b3RE : out sfixed(4 downto -4);
--		b0IM : out sfixed(4 downto -4); 
--		b1IM : out sfixed(4 downto -4); 
--		b2IM : out sfixed(4 downto -4);
--		b3IM : out sfixed(4 downto -4);
		Output: out String(1 to 64);
		finished: out STD_logic:= '0'
	);
end entity;

----------------------------------
--	Architecture Declaration 	--
----------------------------------

architecture compute of qft_2qbit is
 
------------------------
-- signal declaration --
------------------------
type ket is array(0 to 3) of sfixed(4 downto -4);
signal QstateRE, QstateRE_next, QstateIM, QstateIM_next : ket := ("000000000", "000000000", "000000000", "000000000"); -- can this be done in better way ?

type FSM_state_type is (idle,hadamard1,hadamard2,rotation1,swap, Stitch, Convert, finish); -- For 2 qbits 2 hadamard gates and 1 rotation gate.
signal state, state_next : FSM_state_type:=idle;

--type String is array (positive range <>) of character;
signal char0IM, char0RE, char1IM, char1RE, char2IM, char2RE, char3IM, char3RE: String(1 to 8):= "00000000";


------------------------
--      processes     --
------------------------
begin
process(clk,reset)
       begin
            if reset = '0' then
                 state <= idle;
					  --real part
					  QstateRE(0) <= "000010000";--"000011000";--|00> QstateRE(0) = 1.5 in decimal
					  QstateRE(1) <= "000100000";--"000110000";--|01> QstateRE(1) = 3.0 in decimal
					  QstateRE(2) <= "000100000";--"000010100";--|10> QstateRE(2) = 1.25 in decimal
					  QstateRE(3) <= "000110000";--"001000010";--|11> QstateRE(3) = 4.125 in decimal
					  --imaginary part
					  QstateIM(0) <= "000110000";--"000010001";--|00> QstateIM(0) = 1.0625 in decimal
					  QstateIM(1) <= "000010000";--"000100010";--|01> QstateIM(1) = 2.125 in decimal
					  QstateIM(2) <= "000100000";--"000001000";--|10> QstateIM(2) = 0.5 in decimal
					  QstateIM(3) <= "000010000";--"001010000";--|11> QstateIM(3) = 5.0 in decimal
           elsif clk = '1' and clk'event then --falling_edge(clk) then --
                 state<=state_next;
					  QstateRE <= QstateRE_next;
					  QstateIM <= QstateIM_next;
           end if;
       end process;
 
	QFT : process( clk, state, start )
	variable temp1RE,temp2RE,temp3RE,temp4RE : sfixed(5 downto -4) := "0000000000";
	variable temp1IM,temp2IM,temp3IM,temp4IM : sfixed(5 downto -4) := "0000000000";
	begin
	-- avoid latch ( I'm not sure why this is done)
      state_next<=state;
		QstateRE_next<=QstateRE;
		QstateIM_next<=QstateIM;
	--FSM
		case state is
		when idle =>
			if start ='0' then
				state_next <= hadamard1;
			else 
				state_next <= idle;
			end if;
		when hadamard1 =>
			 --calculate real part
			 temp1RE := QstateRE(0) + QstateRE(2);
			 temp2RE := QstateRE(1) + QstateRE(3);
			 temp3RE := QstateRE(0) - QstateRE(2);
			 temp4RE := QstateRE(1) - QstateRE(3);			 
			 --calculate imagniary part
			 temp1IM := QstateIM(0) + QstateIM(2);
			 temp2IM := QstateIM(1) + QstateIM(3);
			 temp3IM := QstateIM(0) - QstateIM(2);
			 temp4IM := QstateIM(1) - QstateIM(3);		 
			 --update ket
			 QstateRE_next(0) <= resize(temp1RE,QstateRE_next(0));--temp1RE(4 downto -4);
			 QstateRE_next(1) <= resize(temp2RE,QstateRE_next(1));--temp2RE(4 downto -4);
			 QstateRE_next(2) <= resize(temp3RE,QstateRE_next(2));--temp3RE(4 downto -4);
			 QstateRE_next(3) <= resize(temp4RE,QstateRE_next(3));--temp4RE(4 downto -4);
			 
			 QstateIM_next(0) <= resize(temp1IM,QstateIM_next(0));--temp1IM(4 downto -4);
			 QstateIM_next(1) <= resize(temp2IM,QstateIM_next(1));--temp2IM(4 downto -4);
			 QstateIM_next(2) <= resize(temp3IM,QstateIM_next(2));--temp3IM(4 downto -4);
			 QstateIM_next(3) <= resize(temp4IM,QstateIM_next(3));--temp4IM(4 downto -4);
			 
			 --next state
			 state_next <= rotation1;
			 
			 
		when rotation1 =>
			 --calculate
			 temp4RE := -QstateIM(3);
			 --update ket
			 QstateRE_next(3) <= resize(temp4RE,QstateRE_next(3));
			 QstateIM_next(3) <= QstateRE(3);
			 --next state
			 state_next <= hadamard2;
			 
		when hadamard2 =>
			 --calculate real part		
			 temp1RE := QstateRE(0) + QstateRE(1);
			 temp2RE := QstateRE(0) - QstateRE(1);
			 temp3RE := QstateRE(2) + QstateRE(3);
			 temp4RE := QstateRE(2) - QstateRE(3);
			 --calculate imagniary part
			 temp1IM := QstateIM(0) + QstateIM(1);
			 temp2IM := QstateIM(0) - QstateIM(1);
			 temp3IM := QstateIM(2) + QstateIM(3);
			 temp4IM := QstateIM(2) - QstateIM(3);	
			 --update ket
			 QstateRE_next(0) <= resize(temp1RE,QstateRE_next(0));--temp1RE(4 downto -4);
			 QstateRE_next(1) <= resize(temp2RE,QstateRE_next(1));--temp2RE(4 downto -4);
			 QstateRE_next(2) <= resize(temp3RE,QstateRE_next(2));--temp3RE(4 downto -4);
			 QstateRE_next(3) <= resize(temp4RE,QstateRE_next(3));--temp4RE(4 downto -4);
			 
			 QstateIM_next(0) <= resize(temp1IM,QstateIM_next(0));--temp1IM(4 downto -4);
			 QstateIM_next(1) <= resize(temp2IM,QstateIM_next(1));--temp2IM(4 downto -4);
			 QstateIM_next(2) <= resize(temp3IM,QstateIM_next(2));--temp3IM(4 downto -4);
			 QstateIM_next(3) <= resize(temp4IM,QstateIM_next(3));--temp4IM(4 downto -4);
			 --next state
			 state_next <= swap;
		
		when swap =>
			QstateRE_next(1) <= QstateRE(2);
			QstateRE_next(2) <= QstateRE(1);
			QstateIM_next(1) <= QstateIM(2);
			QstateIM_next(2) <= QstateIM(1);
			state_next <= Convert;
			 
		when Convert =>
			if QstateRE(0) = to_sfixed(-15.9375,QstateRE(0)) then
				char0RE <= "-15.9375";
			elsif QstateRE(0) = to_sfixed(-15.8750,QstateRE(0)) then
				char0RE <= "-15.8750";
			elsif QstateRE(0) = to_sfixed(-15.8125,QstateRE(0)) then
				char0RE <= "-15.8125";
			elsif QstateRE(0) = to_sfixed(-15.7500,QstateRE(0)) then
				char0RE <= "-15.7500";
			elsif QstateRE(0) = to_sfixed(-15.6875,QstateRE(0)) then
				char0RE <= "-15.6875";
			elsif QstateRE(0) = to_sfixed(-15.6250,QstateRE(0)) then
				char0RE <= "-15.6250";
			elsif QstateRE(0) = to_sfixed(-15.5625,QstateRE(0)) then
				char0RE <= "-15.5625";
			elsif QstateRE(0) = to_sfixed(-15.5000,QstateRE(0)) then
				char0RE <= "-15.5000";
			elsif QstateRE(0) = to_sfixed(-15.4375,QstateRE(0)) then
				char0RE <= "-15.4375";
			elsif QstateRE(0) = to_sfixed(-15.3750,QstateRE(0)) then
				char0RE <= "-15.3750";
			elsif QstateRE(0) = to_sfixed(-15.3125,QstateRE(0)) then
				char0RE <= "-15.3125";
			elsif QstateRE(0) = to_sfixed(-15.2500,QstateRE(0)) then
				char0RE <= "-15.2500";
			elsif QstateRE(0) = to_sfixed(-15.1875,QstateRE(0)) then
				char0RE <= "-15.1875";
			elsif QstateRE(0) = to_sfixed(-15.1250,QstateRE(0)) then
				char0RE <= "-15.1250";
			elsif QstateRE(0) = to_sfixed(-15.0625,QstateRE(0)) then
				char0RE <= "-15.0625";
			elsif QstateRE(0) = to_sfixed(-15.0000,QstateRE(0)) then
				char0RE <= "-15.0000";
			elsif QstateRE(0) = to_sfixed(-14.9375,QstateRE(0)) then
				char0RE <= "-14.9375";
			elsif QstateRE(0) = to_sfixed(-14.8750,QstateRE(0)) then
				char0RE <= "-14.8750";
			elsif QstateRE(0) = to_sfixed(-14.8125,QstateRE(0)) then
				char0RE <= "-14.8125";
			elsif QstateRE(0) = to_sfixed(-14.7500,QstateRE(0)) then
				char0RE <= "-14.7500";
			elsif QstateRE(0) = to_sfixed(-14.6875,QstateRE(0)) then
				char0RE <= "-14.6875";
			elsif QstateRE(0) = to_sfixed(-14.6250,QstateRE(0)) then
				char0RE <= "-14.6250";
			elsif QstateRE(0) = to_sfixed(-14.5625,QstateRE(0)) then
				char0RE <= "-14.5625";
			elsif QstateRE(0) = to_sfixed(-14.5000,QstateRE(0)) then
				char0RE <= "-14.5000";
			elsif QstateRE(0) = to_sfixed(-14.4375,QstateRE(0)) then
				char0RE <= "-14.4375";
			elsif QstateRE(0) = to_sfixed(-14.3750,QstateRE(0)) then
				char0RE <= "-14.3750";
			elsif QstateRE(0) = to_sfixed(-14.3125,QstateRE(0)) then
				char0RE <= "-14.3125";
			elsif QstateRE(0) = to_sfixed(-14.2500,QstateRE(0)) then
				char0RE <= "-14.2500";
			elsif QstateRE(0) = to_sfixed(-14.1875,QstateRE(0)) then
				char0RE <= "-14.1875";
			elsif QstateRE(0) = to_sfixed(-14.1250,QstateRE(0)) then
				char0RE <= "-14.1250";
			elsif QstateRE(0) = to_sfixed(-14.0625,QstateRE(0)) then
				char0RE <= "-14.0625";
			elsif QstateRE(0) = to_sfixed(-14.0000,QstateRE(0)) then
				char0RE <= "-14.0000";
			elsif QstateRE(0) = to_sfixed(-13.9375,QstateRE(0)) then
				char0RE <= "-13.9375";
			elsif QstateRE(0) = to_sfixed(-13.8750,QstateRE(0)) then
				char0RE <= "-13.8750";
			elsif QstateRE(0) = to_sfixed(-13.8125,QstateRE(0)) then
				char0RE <= "-13.8125";
			elsif QstateRE(0) = to_sfixed(-13.7500,QstateRE(0)) then
				char0RE <= "-13.7500";
			elsif QstateRE(0) = to_sfixed(-13.6875,QstateRE(0)) then
				char0RE <= "-13.6875";
			elsif QstateRE(0) = to_sfixed(-13.6250,QstateRE(0)) then
				char0RE <= "-13.6250";
			elsif QstateRE(0) = to_sfixed(-13.5625,QstateRE(0)) then
				char0RE <= "-13.5625";
			elsif QstateRE(0) = to_sfixed(-13.5000,QstateRE(0)) then
				char0RE <= "-13.5000";
			elsif QstateRE(0) = to_sfixed(-13.4375,QstateRE(0)) then
				char0RE <= "-13.4375";
			elsif QstateRE(0) = to_sfixed(-13.3750,QstateRE(0)) then
				char0RE <= "-13.3750";
			elsif QstateRE(0) = to_sfixed(-13.3125,QstateRE(0)) then
				char0RE <= "-13.3125";
			elsif QstateRE(0) = to_sfixed(-13.2500,QstateRE(0)) then
				char0RE <= "-13.2500";
			elsif QstateRE(0) = to_sfixed(-13.1875,QstateRE(0)) then
				char0RE <= "-13.1875";
			elsif QstateRE(0) = to_sfixed(-13.1250,QstateRE(0)) then
				char0RE <= "-13.1250";
			elsif QstateRE(0) = to_sfixed(-13.0625,QstateRE(0)) then
				char0RE <= "-13.0625";
			elsif QstateRE(0) = to_sfixed(-13.0000,QstateRE(0)) then
				char0RE <= "-13.0000";
			elsif QstateRE(0) = to_sfixed(-12.9375,QstateRE(0)) then
				char0RE <= "-12.9375";
			elsif QstateRE(0) = to_sfixed(-12.8750,QstateRE(0)) then
				char0RE <= "-12.8750";
			elsif QstateRE(0) = to_sfixed(-12.8125,QstateRE(0)) then
				char0RE <= "-12.8125";
			elsif QstateRE(0) = to_sfixed(-12.7500,QstateRE(0)) then
				char0RE <= "-12.7500";
			elsif QstateRE(0) = to_sfixed(-12.6875,QstateRE(0)) then
				char0RE <= "-12.6875";
			elsif QstateRE(0) = to_sfixed(-12.6250,QstateRE(0)) then
				char0RE <= "-12.6250";
			elsif QstateRE(0) = to_sfixed(-12.5625,QstateRE(0)) then
				char0RE <= "-12.5625";
			elsif QstateRE(0) = to_sfixed(-12.5000,QstateRE(0)) then
				char0RE <= "-12.5000";
			elsif QstateRE(0) = to_sfixed(-12.4375,QstateRE(0)) then
				char0RE <= "-12.4375";
			elsif QstateRE(0) = to_sfixed(-12.3750,QstateRE(0)) then
				char0RE <= "-12.3750";
			elsif QstateRE(0) = to_sfixed(-12.3125,QstateRE(0)) then
				char0RE <= "-12.3125";
			elsif QstateRE(0) = to_sfixed(-12.2500,QstateRE(0)) then
				char0RE <= "-12.2500";
			elsif QstateRE(0) = to_sfixed(-12.1875,QstateRE(0)) then
				char0RE <= "-12.1875";
			elsif QstateRE(0) = to_sfixed(-12.1250,QstateRE(0)) then
				char0RE <= "-12.1250";
			elsif QstateRE(0) = to_sfixed(-12.0625,QstateRE(0)) then
				char0RE <= "-12.0625";
			elsif QstateRE(0) = to_sfixed(-12.0000,QstateRE(0)) then
				char0RE <= "-12.0000";
			elsif QstateRE(0) = to_sfixed(-11.9375,QstateRE(0)) then
				char0RE <= "-11.9375";
			elsif QstateRE(0) = to_sfixed(-11.8750,QstateRE(0)) then
				char0RE <= "-11.8750";
			elsif QstateRE(0) = to_sfixed(-11.8125,QstateRE(0)) then
				char0RE <= "-11.8125";
			elsif QstateRE(0) = to_sfixed(-11.7500,QstateRE(0)) then
				char0RE <= "-11.7500";
			elsif QstateRE(0) = to_sfixed(-11.6875,QstateRE(0)) then
				char0RE <= "-11.6875";
			elsif QstateRE(0) = to_sfixed(-11.6250,QstateRE(0)) then
				char0RE <= "-11.6250";
			elsif QstateRE(0) = to_sfixed(-11.5625,QstateRE(0)) then
				char0RE <= "-11.5625";
			elsif QstateRE(0) = to_sfixed(-11.5000,QstateRE(0)) then
				char0RE <= "-11.5000";
			elsif QstateRE(0) = to_sfixed(-11.4375,QstateRE(0)) then
				char0RE <= "-11.4375";
			elsif QstateRE(0) = to_sfixed(-11.3750,QstateRE(0)) then
				char0RE <= "-11.3750";
			elsif QstateRE(0) = to_sfixed(-11.3125,QstateRE(0)) then
				char0RE <= "-11.3125";
			elsif QstateRE(0) = to_sfixed(-11.2500,QstateRE(0)) then
				char0RE <= "-11.2500";
			elsif QstateRE(0) = to_sfixed(-11.1875,QstateRE(0)) then
				char0RE <= "-11.1875";
			elsif QstateRE(0) = to_sfixed(-11.1250,QstateRE(0)) then
				char0RE <= "-11.1250";
			elsif QstateRE(0) = to_sfixed(-11.0625,QstateRE(0)) then
				char0RE <= "-11.0625";
			elsif QstateRE(0) = to_sfixed(-11.0000,QstateRE(0)) then
				char0RE <= "-11.0000";
			elsif QstateRE(0) = to_sfixed(-10.9375,QstateRE(0)) then
				char0RE <= "-10.9375";
			elsif QstateRE(0) = to_sfixed(-10.8750,QstateRE(0)) then
				char0RE <= "-10.8750";
			elsif QstateRE(0) = to_sfixed(-10.8125,QstateRE(0)) then
				char0RE <= "-10.8125";
			elsif QstateRE(0) = to_sfixed(-10.7500,QstateRE(0)) then
				char0RE <= "-10.7500";
			elsif QstateRE(0) = to_sfixed(-10.6875,QstateRE(0)) then
				char0RE <= "-10.6875";
			elsif QstateRE(0) = to_sfixed(-10.6250,QstateRE(0)) then
				char0RE <= "-10.6250";
			elsif QstateRE(0) = to_sfixed(-10.5625,QstateRE(0)) then
				char0RE <= "-10.5625";
			elsif QstateRE(0) = to_sfixed(-10.5000,QstateRE(0)) then
				char0RE <= "-10.5000";
			elsif QstateRE(0) = to_sfixed(-10.4375,QstateRE(0)) then
				char0RE <= "-10.4375";
			elsif QstateRE(0) = to_sfixed(-10.3750,QstateRE(0)) then
				char0RE <= "-10.3750";
			elsif QstateRE(0) = to_sfixed(-10.3125,QstateRE(0)) then
				char0RE <= "-10.3125";
			elsif QstateRE(0) = to_sfixed(-10.2500,QstateRE(0)) then
				char0RE <= "-10.2500";
			elsif QstateRE(0) = to_sfixed(-10.1875,QstateRE(0)) then
				char0RE <= "-10.1875";
			elsif QstateRE(0) = to_sfixed(-10.1250,QstateRE(0)) then
				char0RE <= "-10.1250";
			elsif QstateRE(0) = to_sfixed(-10.0625,QstateRE(0)) then
				char0RE <= "-10.0625";
			elsif QstateRE(0) = to_sfixed(-10.0000,QstateRE(0)) then
				char0RE <= "-10.0000";
			elsif QstateRE(0) = to_sfixed(-9.9375,QstateRE(0)) then
				char0RE <= "--9.9375";
			elsif QstateRE(0) = to_sfixed(-9.8750,QstateRE(0)) then
				char0RE <= "--9.8750";
			elsif QstateRE(0) = to_sfixed(-9.8125,QstateRE(0)) then
				char0RE <= "--9.8125";
			elsif QstateRE(0) = to_sfixed(-9.7500,QstateRE(0)) then
				char0RE <= "--9.7500";
			elsif QstateRE(0) = to_sfixed(-9.6875,QstateRE(0)) then
				char0RE <= "--9.6875";
			elsif QstateRE(0) = to_sfixed(-9.6250,QstateRE(0)) then
				char0RE <= "--9.6250";
			elsif QstateRE(0) = to_sfixed(-9.5625,QstateRE(0)) then
				char0RE <= "--9.5625";
			elsif QstateRE(0) = to_sfixed(-9.5000,QstateRE(0)) then
				char0RE <= "--9.5000";
			elsif QstateRE(0) = to_sfixed(-9.4375,QstateRE(0)) then
				char0RE <= "--9.4375";
			elsif QstateRE(0) = to_sfixed(-9.3750,QstateRE(0)) then
				char0RE <= "--9.3750";
			elsif QstateRE(0) = to_sfixed(-9.3125,QstateRE(0)) then
				char0RE <= "--9.3125";
			elsif QstateRE(0) = to_sfixed(-9.2500,QstateRE(0)) then
				char0RE <= "--9.2500";
			elsif QstateRE(0) = to_sfixed(-9.1875,QstateRE(0)) then
				char0RE <= "--9.1875";
			elsif QstateRE(0) = to_sfixed(-9.1250,QstateRE(0)) then
				char0RE <= "--9.1250";
			elsif QstateRE(0) = to_sfixed(-9.0625,QstateRE(0)) then
				char0RE <= "--9.0625";
			elsif QstateRE(0) = to_sfixed(-9.0000,QstateRE(0)) then
				char0RE <= "--9.0000";
			elsif QstateRE(0) = to_sfixed(-8.9375,QstateRE(0)) then
				char0RE <= "--8.9375";
			elsif QstateRE(0) = to_sfixed(-8.8750,QstateRE(0)) then
				char0RE <= "--8.8750";
			elsif QstateRE(0) = to_sfixed(-8.8125,QstateRE(0)) then
				char0RE <= "--8.8125";
			elsif QstateRE(0) = to_sfixed(-8.7500,QstateRE(0)) then
				char0RE <= "--8.7500";
			elsif QstateRE(0) = to_sfixed(-8.6875,QstateRE(0)) then
				char0RE <= "--8.6875";
			elsif QstateRE(0) = to_sfixed(-8.6250,QstateRE(0)) then
				char0RE <= "--8.6250";
			elsif QstateRE(0) = to_sfixed(-8.5625,QstateRE(0)) then
				char0RE <= "--8.5625";
			elsif QstateRE(0) = to_sfixed(-8.5000,QstateRE(0)) then
				char0RE <= "--8.5000";
			elsif QstateRE(0) = to_sfixed(-8.4375,QstateRE(0)) then
				char0RE <= "--8.4375";
			elsif QstateRE(0) = to_sfixed(-8.3750,QstateRE(0)) then
				char0RE <= "--8.3750";
			elsif QstateRE(0) = to_sfixed(-8.3125,QstateRE(0)) then
				char0RE <= "--8.3125";
			elsif QstateRE(0) = to_sfixed(-8.2500,QstateRE(0)) then
				char0RE <= "--8.2500";
			elsif QstateRE(0) = to_sfixed(-8.1875,QstateRE(0)) then
				char0RE <= "--8.1875";
			elsif QstateRE(0) = to_sfixed(-8.1250,QstateRE(0)) then
				char0RE <= "--8.1250";
			elsif QstateRE(0) = to_sfixed(-8.0625,QstateRE(0)) then
				char0RE <= "--8.0625";
			elsif QstateRE(0) = to_sfixed(-8.0000,QstateRE(0)) then
				char0RE <= "--8.0000";
			elsif QstateRE(0) = to_sfixed(-7.9375,QstateRE(0)) then
				char0RE <= "--7.9375";
			elsif QstateRE(0) = to_sfixed(-7.8750,QstateRE(0)) then
				char0RE <= "--7.8750";
			elsif QstateRE(0) = to_sfixed(-7.8125,QstateRE(0)) then
				char0RE <= "--7.8125";
			elsif QstateRE(0) = to_sfixed(-7.7500,QstateRE(0)) then
				char0RE <= "--7.7500";
			elsif QstateRE(0) = to_sfixed(-7.6875,QstateRE(0)) then
				char0RE <= "--7.6875";
			elsif QstateRE(0) = to_sfixed(-7.6250,QstateRE(0)) then
				char0RE <= "--7.6250";
			elsif QstateRE(0) = to_sfixed(-7.5625,QstateRE(0)) then
				char0RE <= "--7.5625";
			elsif QstateRE(0) = to_sfixed(-7.5000,QstateRE(0)) then
				char0RE <= "--7.5000";
			elsif QstateRE(0) = to_sfixed(-7.4375,QstateRE(0)) then
				char0RE <= "--7.4375";
			elsif QstateRE(0) = to_sfixed(-7.3750,QstateRE(0)) then
				char0RE <= "--7.3750";
			elsif QstateRE(0) = to_sfixed(-7.3125,QstateRE(0)) then
				char0RE <= "--7.3125";
			elsif QstateRE(0) = to_sfixed(-7.2500,QstateRE(0)) then
				char0RE <= "--7.2500";
			elsif QstateRE(0) = to_sfixed(-7.1875,QstateRE(0)) then
				char0RE <= "--7.1875";
			elsif QstateRE(0) = to_sfixed(-7.1250,QstateRE(0)) then
				char0RE <= "--7.1250";
			elsif QstateRE(0) = to_sfixed(-7.0625,QstateRE(0)) then
				char0RE <= "--7.0625";
			elsif QstateRE(0) = to_sfixed(-7.0000,QstateRE(0)) then
				char0RE <= "--7.0000";
			elsif QstateRE(0) = to_sfixed(-6.9375,QstateRE(0)) then
				char0RE <= "--6.9375";
			elsif QstateRE(0) = to_sfixed(-6.8750,QstateRE(0)) then
				char0RE <= "--6.8750";
			elsif QstateRE(0) = to_sfixed(-6.8125,QstateRE(0)) then
				char0RE <= "--6.8125";
			elsif QstateRE(0) = to_sfixed(-6.7500,QstateRE(0)) then
				char0RE <= "--6.7500";
			elsif QstateRE(0) = to_sfixed(-6.6875,QstateRE(0)) then
				char0RE <= "--6.6875";
			elsif QstateRE(0) = to_sfixed(-6.6250,QstateRE(0)) then
				char0RE <= "--6.6250";
			elsif QstateRE(0) = to_sfixed(-6.5625,QstateRE(0)) then
				char0RE <= "--6.5625";
			elsif QstateRE(0) = to_sfixed(-6.5000,QstateRE(0)) then
				char0RE <= "--6.5000";
			elsif QstateRE(0) = to_sfixed(-6.4375,QstateRE(0)) then
				char0RE <= "--6.4375";
			elsif QstateRE(0) = to_sfixed(-6.3750,QstateRE(0)) then
				char0RE <= "--6.3750";
			elsif QstateRE(0) = to_sfixed(-6.3125,QstateRE(0)) then
				char0RE <= "--6.3125";
			elsif QstateRE(0) = to_sfixed(-6.2500,QstateRE(0)) then
				char0RE <= "--6.2500";
			elsif QstateRE(0) = to_sfixed(-6.1875,QstateRE(0)) then
				char0RE <= "--6.1875";
			elsif QstateRE(0) = to_sfixed(-6.1250,QstateRE(0)) then
				char0RE <= "--6.1250";
			elsif QstateRE(0) = to_sfixed(-6.0625,QstateRE(0)) then
				char0RE <= "--6.0625";
			elsif QstateRE(0) = to_sfixed(-6.0000,QstateRE(0)) then
				char0RE <= "--6.0000";
			elsif QstateRE(0) = to_sfixed(-5.9375,QstateRE(0)) then
				char0RE <= "--5.9375";
			elsif QstateRE(0) = to_sfixed(-5.8750,QstateRE(0)) then
				char0RE <= "--5.8750";
			elsif QstateRE(0) = to_sfixed(-5.8125,QstateRE(0)) then
				char0RE <= "--5.8125";
			elsif QstateRE(0) = to_sfixed(-5.7500,QstateRE(0)) then
				char0RE <= "--5.7500";
			elsif QstateRE(0) = to_sfixed(-5.6875,QstateRE(0)) then
				char0RE <= "--5.6875";
			elsif QstateRE(0) = to_sfixed(-5.6250,QstateRE(0)) then
				char0RE <= "--5.6250";
			elsif QstateRE(0) = to_sfixed(-5.5625,QstateRE(0)) then
				char0RE <= "--5.5625";
			elsif QstateRE(0) = to_sfixed(-5.5000,QstateRE(0)) then
				char0RE <= "--5.5000";
			elsif QstateRE(0) = to_sfixed(-5.4375,QstateRE(0)) then
				char0RE <= "--5.4375";
			elsif QstateRE(0) = to_sfixed(-5.3750,QstateRE(0)) then
				char0RE <= "--5.3750";
			elsif QstateRE(0) = to_sfixed(-5.3125,QstateRE(0)) then
				char0RE <= "--5.3125";
			elsif QstateRE(0) = to_sfixed(-5.2500,QstateRE(0)) then
				char0RE <= "--5.2500";
			elsif QstateRE(0) = to_sfixed(-5.1875,QstateRE(0)) then
				char0RE <= "--5.1875";
			elsif QstateRE(0) = to_sfixed(-5.1250,QstateRE(0)) then
				char0RE <= "--5.1250";
			elsif QstateRE(0) = to_sfixed(-5.0625,QstateRE(0)) then
				char0RE <= "--5.0625";
			elsif QstateRE(0) = to_sfixed(-5.0000,QstateRE(0)) then
				char0RE <= "--5.0000";
			elsif QstateRE(0) = to_sfixed(-4.9375,QstateRE(0)) then
				char0RE <= "--4.9375";
			elsif QstateRE(0) = to_sfixed(-4.8750,QstateRE(0)) then
				char0RE <= "--4.8750";
			elsif QstateRE(0) = to_sfixed(-4.8125,QstateRE(0)) then
				char0RE <= "--4.8125";
			elsif QstateRE(0) = to_sfixed(-4.7500,QstateRE(0)) then
				char0RE <= "--4.7500";
			elsif QstateRE(0) = to_sfixed(-4.6875,QstateRE(0)) then
				char0RE <= "--4.6875";
			elsif QstateRE(0) = to_sfixed(-4.6250,QstateRE(0)) then
				char0RE <= "--4.6250";
			elsif QstateRE(0) = to_sfixed(-4.5625,QstateRE(0)) then
				char0RE <= "--4.5625";
			elsif QstateRE(0) = to_sfixed(-4.5000,QstateRE(0)) then
				char0RE <= "--4.5000";
			elsif QstateRE(0) = to_sfixed(-4.4375,QstateRE(0)) then
				char0RE <= "--4.4375";
			elsif QstateRE(0) = to_sfixed(-4.3750,QstateRE(0)) then
				char0RE <= "--4.3750";
			elsif QstateRE(0) = to_sfixed(-4.3125,QstateRE(0)) then
				char0RE <= "--4.3125";
			elsif QstateRE(0) = to_sfixed(-4.2500,QstateRE(0)) then
				char0RE <= "--4.2500";
			elsif QstateRE(0) = to_sfixed(-4.1875,QstateRE(0)) then
				char0RE <= "--4.1875";
			elsif QstateRE(0) = to_sfixed(-4.1250,QstateRE(0)) then
				char0RE <= "--4.1250";
			elsif QstateRE(0) = to_sfixed(-4.0625,QstateRE(0)) then
				char0RE <= "--4.0625";
			elsif QstateRE(0) = to_sfixed(-4.0000,QstateRE(0)) then
				char0RE <= "--4.0000";
			elsif QstateRE(0) = to_sfixed(-3.9375,QstateRE(0)) then
				char0RE <= "--3.9375";
			elsif QstateRE(0) = to_sfixed(-3.8750,QstateRE(0)) then
				char0RE <= "--3.8750";
			elsif QstateRE(0) = to_sfixed(-3.8125,QstateRE(0)) then
				char0RE <= "--3.8125";
			elsif QstateRE(0) = to_sfixed(-3.7500,QstateRE(0)) then
				char0RE <= "--3.7500";
			elsif QstateRE(0) = to_sfixed(-3.6875,QstateRE(0)) then
				char0RE <= "--3.6875";
			elsif QstateRE(0) = to_sfixed(-3.6250,QstateRE(0)) then
				char0RE <= "--3.6250";
			elsif QstateRE(0) = to_sfixed(-3.5625,QstateRE(0)) then
				char0RE <= "--3.5625";
			elsif QstateRE(0) = to_sfixed(-3.5000,QstateRE(0)) then
				char0RE <= "--3.5000";
			elsif QstateRE(0) = to_sfixed(-3.4375,QstateRE(0)) then
				char0RE <= "--3.4375";
			elsif QstateRE(0) = to_sfixed(-3.3750,QstateRE(0)) then
				char0RE <= "--3.3750";
			elsif QstateRE(0) = to_sfixed(-3.3125,QstateRE(0)) then
				char0RE <= "--3.3125";
			elsif QstateRE(0) = to_sfixed(-3.2500,QstateRE(0)) then
				char0RE <= "--3.2500";
			elsif QstateRE(0) = to_sfixed(-3.1875,QstateRE(0)) then
				char0RE <= "--3.1875";
			elsif QstateRE(0) = to_sfixed(-3.1250,QstateRE(0)) then
				char0RE <= "--3.1250";
			elsif QstateRE(0) = to_sfixed(-3.0625,QstateRE(0)) then
				char0RE <= "--3.0625";
			elsif QstateRE(0) = to_sfixed(-3.0000,QstateRE(0)) then
				char0RE <= "--3.0000";
			elsif QstateRE(0) = to_sfixed(-2.9375,QstateRE(0)) then
				char0RE <= "--2.9375";
			elsif QstateRE(0) = to_sfixed(-2.8750,QstateRE(0)) then
				char0RE <= "--2.8750";
			elsif QstateRE(0) = to_sfixed(-2.8125,QstateRE(0)) then
				char0RE <= "--2.8125";
			elsif QstateRE(0) = to_sfixed(-2.7500,QstateRE(0)) then
				char0RE <= "--2.7500";
			elsif QstateRE(0) = to_sfixed(-2.6875,QstateRE(0)) then
				char0RE <= "--2.6875";
			elsif QstateRE(0) = to_sfixed(-2.6250,QstateRE(0)) then
				char0RE <= "--2.6250";
			elsif QstateRE(0) = to_sfixed(-2.5625,QstateRE(0)) then
				char0RE <= "--2.5625";
			elsif QstateRE(0) = to_sfixed(-2.5000,QstateRE(0)) then
				char0RE <= "--2.5000";
			elsif QstateRE(0) = to_sfixed(-2.4375,QstateRE(0)) then
				char0RE <= "--2.4375";
			elsif QstateRE(0) = to_sfixed(-2.3750,QstateRE(0)) then
				char0RE <= "--2.3750";
			elsif QstateRE(0) = to_sfixed(-2.3125,QstateRE(0)) then
				char0RE <= "--2.3125";
			elsif QstateRE(0) = to_sfixed(-2.2500,QstateRE(0)) then
				char0RE <= "--2.2500";
			elsif QstateRE(0) = to_sfixed(-2.1875,QstateRE(0)) then
				char0RE <= "--2.1875";
			elsif QstateRE(0) = to_sfixed(-2.1250,QstateRE(0)) then
				char0RE <= "--2.1250";
			elsif QstateRE(0) = to_sfixed(-2.0625,QstateRE(0)) then
				char0RE <= "--2.0625";
			elsif QstateRE(0) = to_sfixed(-2.0000,QstateRE(0)) then
				char0RE <= "--2.0000";
			elsif QstateRE(0) = to_sfixed(-1.9375,QstateRE(0)) then
				char0RE <= "--1.9375";
			elsif QstateRE(0) = to_sfixed(-1.8750,QstateRE(0)) then
				char0RE <= "--1.8750";
			elsif QstateRE(0) = to_sfixed(-1.8125,QstateRE(0)) then
				char0RE <= "--1.8125";
			elsif QstateRE(0) = to_sfixed(-1.7500,QstateRE(0)) then
				char0RE <= "--1.7500";
			elsif QstateRE(0) = to_sfixed(-1.6875,QstateRE(0)) then
				char0RE <= "--1.6875";
			elsif QstateRE(0) = to_sfixed(-1.6250,QstateRE(0)) then
				char0RE <= "--1.6250";
			elsif QstateRE(0) = to_sfixed(-1.5625,QstateRE(0)) then
				char0RE <= "--1.5625";
			elsif QstateRE(0) = to_sfixed(-1.5000,QstateRE(0)) then
				char0RE <= "--1.5000";
			elsif QstateRE(0) = to_sfixed(-1.4375,QstateRE(0)) then
				char0RE <= "--1.4375";
			elsif QstateRE(0) = to_sfixed(-1.3750,QstateRE(0)) then
				char0RE <= "--1.3750";
			elsif QstateRE(0) = to_sfixed(-1.3125,QstateRE(0)) then
				char0RE <= "--1.3125";
			elsif QstateRE(0) = to_sfixed(-1.2500,QstateRE(0)) then
				char0RE <= "--1.2500";
			elsif QstateRE(0) = to_sfixed(-1.1875,QstateRE(0)) then
				char0RE <= "--1.1875";
			elsif QstateRE(0) = to_sfixed(-1.1250,QstateRE(0)) then
				char0RE <= "--1.1250";
			elsif QstateRE(0) = to_sfixed(-1.0625,QstateRE(0)) then
				char0RE <= "--1.0625";
			elsif QstateRE(0) = to_sfixed(-1.0000,QstateRE(0)) then
				char0RE <= "--1.0000";
			elsif QstateRE(0) = to_sfixed(-0.9375,QstateRE(0)) then
				char0RE <= "--0.9375";
			elsif QstateRE(0) = to_sfixed(-0.8750,QstateRE(0)) then
				char0RE <= "--0.8750";
			elsif QstateRE(0) = to_sfixed(-0.8125,QstateRE(0)) then
				char0RE <= "--0.8125";
			elsif QstateRE(0) = to_sfixed(-0.7500,QstateRE(0)) then
				char0RE <= "--0.7500";
			elsif QstateRE(0) = to_sfixed(-0.6875,QstateRE(0)) then
				char0RE <= "--0.6875";
			elsif QstateRE(0) = to_sfixed(-0.6250,QstateRE(0)) then
				char0RE <= "--0.6250";
			elsif QstateRE(0) = to_sfixed(-0.5625,QstateRE(0)) then
				char0RE <= "--0.5625";
			elsif QstateRE(0) = to_sfixed(-0.5000,QstateRE(0)) then
				char0RE <= "--0.5000";
			elsif QstateRE(0) = to_sfixed(-0.4375,QstateRE(0)) then
				char0RE <= "--0.4375";
			elsif QstateRE(0) = to_sfixed(-0.3750,QstateRE(0)) then
				char0RE <= "--0.3750";
			elsif QstateRE(0) = to_sfixed(-0.3125,QstateRE(0)) then
				char0RE <= "--0.3125";
			elsif QstateRE(0) = to_sfixed(-0.2500,QstateRE(0)) then
				char0RE <= "--0.2500";
			elsif QstateRE(0) = to_sfixed(-0.1875,QstateRE(0)) then
				char0RE <= "--0.1875";
			elsif QstateRE(0) = to_sfixed(-0.1250,QstateRE(0)) then
				char0RE <= "--0.1250";
			elsif QstateRE(0) = to_sfixed(-0.0625,QstateRE(0)) then
				char0RE <= "--0.0625";
			elsif QstateRE(0) = to_sfixed(00.0000,QstateRE(0)) then
				char0RE <= "+00.0000";
			elsif QstateRE(0) = to_sfixed(00.0625,QstateRE(0)) then
				char0RE <= "+00.0625";
			elsif QstateRE(0) = to_sfixed(00.1250,QstateRE(0)) then
				char0RE <= "+00.1250";
			elsif QstateRE(0) = to_sfixed(00.1875,QstateRE(0)) then
				char0RE <= "+00.1875";
			elsif QstateRE(0) = to_sfixed(00.2500,QstateRE(0)) then
				char0RE <= "+00.2500";
			elsif QstateRE(0) = to_sfixed(00.3125,QstateRE(0)) then
				char0RE <= "+00.3125";
			elsif QstateRE(0) = to_sfixed(00.3750,QstateRE(0)) then
				char0RE <= "+00.3750";
			elsif QstateRE(0) = to_sfixed(00.4375,QstateRE(0)) then
				char0RE <= "+00.4375";
			elsif QstateRE(0) = to_sfixed(00.5000,QstateRE(0)) then
				char0RE <= "+00.5000";
			elsif QstateRE(0) = to_sfixed(00.5625,QstateRE(0)) then
				char0RE <= "+00.5625";
			elsif QstateRE(0) = to_sfixed(00.6250,QstateRE(0)) then
				char0RE <= "+00.6250";
			elsif QstateRE(0) = to_sfixed(00.6875,QstateRE(0)) then
				char0RE <= "+00.6875";
			elsif QstateRE(0) = to_sfixed(00.7500,QstateRE(0)) then
				char0RE <= "+00.7500";
			elsif QstateRE(0) = to_sfixed(00.8125,QstateRE(0)) then
				char0RE <= "+00.8125";
			elsif QstateRE(0) = to_sfixed(00.8750,QstateRE(0)) then
				char0RE <= "+00.8750";
			elsif QstateRE(0) = to_sfixed(00.9375,QstateRE(0)) then
				char0RE <= "+00.9375";
			elsif QstateRE(0) = to_sfixed(01.0000,QstateRE(0)) then
				char0RE <= "+01.0000";
			elsif QstateRE(0) = to_sfixed(01.0625,QstateRE(0)) then
				char0RE <= "+01.0625";
			elsif QstateRE(0) = to_sfixed(01.1250,QstateRE(0)) then
				char0RE <= "+01.1250";
			elsif QstateRE(0) = to_sfixed(01.1875,QstateRE(0)) then
				char0RE <= "+01.1875";
			elsif QstateRE(0) = to_sfixed(01.2500,QstateRE(0)) then
				char0RE <= "+01.2500";
			elsif QstateRE(0) = to_sfixed(01.3125,QstateRE(0)) then
				char0RE <= "+01.3125";
			elsif QstateRE(0) = to_sfixed(01.3750,QstateRE(0)) then
				char0RE <= "+01.3750";
			elsif QstateRE(0) = to_sfixed(01.4375,QstateRE(0)) then
				char0RE <= "+01.4375";
			elsif QstateRE(0) = to_sfixed(01.5000,QstateRE(0)) then
				char0RE <= "+01.5000";
			elsif QstateRE(0) = to_sfixed(01.5625,QstateRE(0)) then
				char0RE <= "+01.5625";
			elsif QstateRE(0) = to_sfixed(01.6250,QstateRE(0)) then
				char0RE <= "+01.6250";
			elsif QstateRE(0) = to_sfixed(01.6875,QstateRE(0)) then
				char0RE <= "+01.6875";
			elsif QstateRE(0) = to_sfixed(01.7500,QstateRE(0)) then
				char0RE <= "+01.7500";
			elsif QstateRE(0) = to_sfixed(01.8125,QstateRE(0)) then
				char0RE <= "+01.8125";
			elsif QstateRE(0) = to_sfixed(01.8750,QstateRE(0)) then
				char0RE <= "+01.8750";
			elsif QstateRE(0) = to_sfixed(01.9375,QstateRE(0)) then
				char0RE <= "+01.9375";
			elsif QstateRE(0) = to_sfixed(02.0000,QstateRE(0)) then
				char0RE <= "+02.0000";
			elsif QstateRE(0) = to_sfixed(02.0625,QstateRE(0)) then
				char0RE <= "+02.0625";
			elsif QstateRE(0) = to_sfixed(02.1250,QstateRE(0)) then
				char0RE <= "+02.1250";
			elsif QstateRE(0) = to_sfixed(02.1875,QstateRE(0)) then
				char0RE <= "+02.1875";
			elsif QstateRE(0) = to_sfixed(02.2500,QstateRE(0)) then
				char0RE <= "+02.2500";
			elsif QstateRE(0) = to_sfixed(02.3125,QstateRE(0)) then
				char0RE <= "+02.3125";
			elsif QstateRE(0) = to_sfixed(02.3750,QstateRE(0)) then
				char0RE <= "+02.3750";
			elsif QstateRE(0) = to_sfixed(02.4375,QstateRE(0)) then
				char0RE <= "+02.4375";
			elsif QstateRE(0) = to_sfixed(02.5000,QstateRE(0)) then
				char0RE <= "+02.5000";
			elsif QstateRE(0) = to_sfixed(02.5625,QstateRE(0)) then
				char0RE <= "+02.5625";
			elsif QstateRE(0) = to_sfixed(02.6250,QstateRE(0)) then
				char0RE <= "+02.6250";
			elsif QstateRE(0) = to_sfixed(02.6875,QstateRE(0)) then
				char0RE <= "+02.6875";
			elsif QstateRE(0) = to_sfixed(02.7500,QstateRE(0)) then
				char0RE <= "+02.7500";
			elsif QstateRE(0) = to_sfixed(02.8125,QstateRE(0)) then
				char0RE <= "+02.8125";
			elsif QstateRE(0) = to_sfixed(02.8750,QstateRE(0)) then
				char0RE <= "+02.8750";
			elsif QstateRE(0) = to_sfixed(02.9375,QstateRE(0)) then
				char0RE <= "+02.9375";
			elsif QstateRE(0) = to_sfixed(03.0000,QstateRE(0)) then
				char0RE <= "+03.0000";
			elsif QstateRE(0) = to_sfixed(03.0625,QstateRE(0)) then
				char0RE <= "+03.0625";
			elsif QstateRE(0) = to_sfixed(03.1250,QstateRE(0)) then
				char0RE <= "+03.1250";
			elsif QstateRE(0) = to_sfixed(03.1875,QstateRE(0)) then
				char0RE <= "+03.1875";
			elsif QstateRE(0) = to_sfixed(03.2500,QstateRE(0)) then
				char0RE <= "+03.2500";
			elsif QstateRE(0) = to_sfixed(03.3125,QstateRE(0)) then
				char0RE <= "+03.3125";
			elsif QstateRE(0) = to_sfixed(03.3750,QstateRE(0)) then
				char0RE <= "+03.3750";
			elsif QstateRE(0) = to_sfixed(03.4375,QstateRE(0)) then
				char0RE <= "+03.4375";
			elsif QstateRE(0) = to_sfixed(03.5000,QstateRE(0)) then
				char0RE <= "+03.5000";
			elsif QstateRE(0) = to_sfixed(03.5625,QstateRE(0)) then
				char0RE <= "+03.5625";
			elsif QstateRE(0) = to_sfixed(03.6250,QstateRE(0)) then
				char0RE <= "+03.6250";
			elsif QstateRE(0) = to_sfixed(03.6875,QstateRE(0)) then
				char0RE <= "+03.6875";
			elsif QstateRE(0) = to_sfixed(03.7500,QstateRE(0)) then
				char0RE <= "+03.7500";
			elsif QstateRE(0) = to_sfixed(03.8125,QstateRE(0)) then
				char0RE <= "+03.8125";
			elsif QstateRE(0) = to_sfixed(03.8750,QstateRE(0)) then
				char0RE <= "+03.8750";
			elsif QstateRE(0) = to_sfixed(03.9375,QstateRE(0)) then
				char0RE <= "+03.9375";
			elsif QstateRE(0) = to_sfixed(04.0000,QstateRE(0)) then
				char0RE <= "+04.0000";
			elsif QstateRE(0) = to_sfixed(04.0625,QstateRE(0)) then
				char0RE <= "+04.0625";
			elsif QstateRE(0) = to_sfixed(04.1250,QstateRE(0)) then
				char0RE <= "+04.1250";
			elsif QstateRE(0) = to_sfixed(04.1875,QstateRE(0)) then
				char0RE <= "+04.1875";
			elsif QstateRE(0) = to_sfixed(04.2500,QstateRE(0)) then
				char0RE <= "+04.2500";
			elsif QstateRE(0) = to_sfixed(04.3125,QstateRE(0)) then
				char0RE <= "+04.3125";
			elsif QstateRE(0) = to_sfixed(04.3750,QstateRE(0)) then
				char0RE <= "+04.3750";
			elsif QstateRE(0) = to_sfixed(04.4375,QstateRE(0)) then
				char0RE <= "+04.4375";
			elsif QstateRE(0) = to_sfixed(04.5000,QstateRE(0)) then
				char0RE <= "+04.5000";
			elsif QstateRE(0) = to_sfixed(04.5625,QstateRE(0)) then
				char0RE <= "+04.5625";
			elsif QstateRE(0) = to_sfixed(04.6250,QstateRE(0)) then
				char0RE <= "+04.6250";
			elsif QstateRE(0) = to_sfixed(04.6875,QstateRE(0)) then
				char0RE <= "+04.6875";
			elsif QstateRE(0) = to_sfixed(04.7500,QstateRE(0)) then
				char0RE <= "+04.7500";
			elsif QstateRE(0) = to_sfixed(04.8125,QstateRE(0)) then
				char0RE <= "+04.8125";
			elsif QstateRE(0) = to_sfixed(04.8750,QstateRE(0)) then
				char0RE <= "+04.8750";
			elsif QstateRE(0) = to_sfixed(04.9375,QstateRE(0)) then
				char0RE <= "+04.9375";
			elsif QstateRE(0) = to_sfixed(05.0000,QstateRE(0)) then
				char0RE <= "+05.0000";
			elsif QstateRE(0) = to_sfixed(05.0625,QstateRE(0)) then
				char0RE <= "+05.0625";
			elsif QstateRE(0) = to_sfixed(05.1250,QstateRE(0)) then
				char0RE <= "+05.1250";
			elsif QstateRE(0) = to_sfixed(05.1875,QstateRE(0)) then
				char0RE <= "+05.1875";
			elsif QstateRE(0) = to_sfixed(05.2500,QstateRE(0)) then
				char0RE <= "+05.2500";
			elsif QstateRE(0) = to_sfixed(05.3125,QstateRE(0)) then
				char0RE <= "+05.3125";
			elsif QstateRE(0) = to_sfixed(05.3750,QstateRE(0)) then
				char0RE <= "+05.3750";
			elsif QstateRE(0) = to_sfixed(05.4375,QstateRE(0)) then
				char0RE <= "+05.4375";
			elsif QstateRE(0) = to_sfixed(05.5000,QstateRE(0)) then
				char0RE <= "+05.5000";
			elsif QstateRE(0) = to_sfixed(05.5625,QstateRE(0)) then
				char0RE <= "+05.5625";
			elsif QstateRE(0) = to_sfixed(05.6250,QstateRE(0)) then
				char0RE <= "+05.6250";
			elsif QstateRE(0) = to_sfixed(05.6875,QstateRE(0)) then
				char0RE <= "+05.6875";
			elsif QstateRE(0) = to_sfixed(05.7500,QstateRE(0)) then
				char0RE <= "+05.7500";
			elsif QstateRE(0) = to_sfixed(05.8125,QstateRE(0)) then
				char0RE <= "+05.8125";
			elsif QstateRE(0) = to_sfixed(05.8750,QstateRE(0)) then
				char0RE <= "+05.8750";
			elsif QstateRE(0) = to_sfixed(05.9375,QstateRE(0)) then
				char0RE <= "+05.9375";
			elsif QstateRE(0) = to_sfixed(06.0000,QstateRE(0)) then
				char0RE <= "+06.0000";
			elsif QstateRE(0) = to_sfixed(06.0625,QstateRE(0)) then
				char0RE <= "+06.0625";
			elsif QstateRE(0) = to_sfixed(06.1250,QstateRE(0)) then
				char0RE <= "+06.1250";
			elsif QstateRE(0) = to_sfixed(06.1875,QstateRE(0)) then
				char0RE <= "+06.1875";
			elsif QstateRE(0) = to_sfixed(06.2500,QstateRE(0)) then
				char0RE <= "+06.2500";
			elsif QstateRE(0) = to_sfixed(06.3125,QstateRE(0)) then
				char0RE <= "+06.3125";
			elsif QstateRE(0) = to_sfixed(06.3750,QstateRE(0)) then
				char0RE <= "+06.3750";
			elsif QstateRE(0) = to_sfixed(06.4375,QstateRE(0)) then
				char0RE <= "+06.4375";
			elsif QstateRE(0) = to_sfixed(06.5000,QstateRE(0)) then
				char0RE <= "+06.5000";
			elsif QstateRE(0) = to_sfixed(06.5625,QstateRE(0)) then
				char0RE <= "+06.5625";
			elsif QstateRE(0) = to_sfixed(06.6250,QstateRE(0)) then
				char0RE <= "+06.6250";
			elsif QstateRE(0) = to_sfixed(06.6875,QstateRE(0)) then
				char0RE <= "+06.6875";
			elsif QstateRE(0) = to_sfixed(06.7500,QstateRE(0)) then
				char0RE <= "+06.7500";
			elsif QstateRE(0) = to_sfixed(06.8125,QstateRE(0)) then
				char0RE <= "+06.8125";
			elsif QstateRE(0) = to_sfixed(06.8750,QstateRE(0)) then
				char0RE <= "+06.8750";
			elsif QstateRE(0) = to_sfixed(06.9375,QstateRE(0)) then
				char0RE <= "+06.9375";
			elsif QstateRE(0) = to_sfixed(07.0000,QstateRE(0)) then
				char0RE <= "+07.0000";
			elsif QstateRE(0) = to_sfixed(07.0625,QstateRE(0)) then
				char0RE <= "+07.0625";
			elsif QstateRE(0) = to_sfixed(07.1250,QstateRE(0)) then
				char0RE <= "+07.1250";
			elsif QstateRE(0) = to_sfixed(07.1875,QstateRE(0)) then
				char0RE <= "+07.1875";
			elsif QstateRE(0) = to_sfixed(07.2500,QstateRE(0)) then
				char0RE <= "+07.2500";
			elsif QstateRE(0) = to_sfixed(07.3125,QstateRE(0)) then
				char0RE <= "+07.3125";
			elsif QstateRE(0) = to_sfixed(07.3750,QstateRE(0)) then
				char0RE <= "+07.3750";
			elsif QstateRE(0) = to_sfixed(07.4375,QstateRE(0)) then
				char0RE <= "+07.4375";
			elsif QstateRE(0) = to_sfixed(07.5000,QstateRE(0)) then
				char0RE <= "+07.5000";
			elsif QstateRE(0) = to_sfixed(07.5625,QstateRE(0)) then
				char0RE <= "+07.5625";
			elsif QstateRE(0) = to_sfixed(07.6250,QstateRE(0)) then
				char0RE <= "+07.6250";
			elsif QstateRE(0) = to_sfixed(07.6875,QstateRE(0)) then
				char0RE <= "+07.6875";
			elsif QstateRE(0) = to_sfixed(07.7500,QstateRE(0)) then
				char0RE <= "+07.7500";
			elsif QstateRE(0) = to_sfixed(07.8125,QstateRE(0)) then
				char0RE <= "+07.8125";
			elsif QstateRE(0) = to_sfixed(07.8750,QstateRE(0)) then
				char0RE <= "+07.8750";
			elsif QstateRE(0) = to_sfixed(07.9375,QstateRE(0)) then
				char0RE <= "+07.9375";
			elsif QstateRE(0) = to_sfixed(08.0000,QstateRE(0)) then
				char0RE <= "+08.0000";
			elsif QstateRE(0) = to_sfixed(08.0625,QstateRE(0)) then
				char0RE <= "+08.0625";
			elsif QstateRE(0) = to_sfixed(08.1250,QstateRE(0)) then
				char0RE <= "+08.1250";
			elsif QstateRE(0) = to_sfixed(08.1875,QstateRE(0)) then
				char0RE <= "+08.1875";
			elsif QstateRE(0) = to_sfixed(08.2500,QstateRE(0)) then
				char0RE <= "+08.2500";
			elsif QstateRE(0) = to_sfixed(08.3125,QstateRE(0)) then
				char0RE <= "+08.3125";
			elsif QstateRE(0) = to_sfixed(08.3750,QstateRE(0)) then
				char0RE <= "+08.3750";
			elsif QstateRE(0) = to_sfixed(08.4375,QstateRE(0)) then
				char0RE <= "+08.4375";
			elsif QstateRE(0) = to_sfixed(08.5000,QstateRE(0)) then
				char0RE <= "+08.5000";
			elsif QstateRE(0) = to_sfixed(08.5625,QstateRE(0)) then
				char0RE <= "+08.5625";
			elsif QstateRE(0) = to_sfixed(08.6250,QstateRE(0)) then
				char0RE <= "+08.6250";
			elsif QstateRE(0) = to_sfixed(08.6875,QstateRE(0)) then
				char0RE <= "+08.6875";
			elsif QstateRE(0) = to_sfixed(08.7500,QstateRE(0)) then
				char0RE <= "+08.7500";
			elsif QstateRE(0) = to_sfixed(08.8125,QstateRE(0)) then
				char0RE <= "+08.8125";
			elsif QstateRE(0) = to_sfixed(08.8750,QstateRE(0)) then
				char0RE <= "+08.8750";
			elsif QstateRE(0) = to_sfixed(08.9375,QstateRE(0)) then
				char0RE <= "+08.9375";
			elsif QstateRE(0) = to_sfixed(09.0000,QstateRE(0)) then
				char0RE <= "+09.0000";
			elsif QstateRE(0) = to_sfixed(09.0625,QstateRE(0)) then
				char0RE <= "+09.0625";
			elsif QstateRE(0) = to_sfixed(09.1250,QstateRE(0)) then
				char0RE <= "+09.1250";
			elsif QstateRE(0) = to_sfixed(09.1875,QstateRE(0)) then
				char0RE <= "+09.1875";
			elsif QstateRE(0) = to_sfixed(09.2500,QstateRE(0)) then
				char0RE <= "+09.2500";
			elsif QstateRE(0) = to_sfixed(09.3125,QstateRE(0)) then
				char0RE <= "+09.3125";
			elsif QstateRE(0) = to_sfixed(09.3750,QstateRE(0)) then
				char0RE <= "+09.3750";
			elsif QstateRE(0) = to_sfixed(09.4375,QstateRE(0)) then
				char0RE <= "+09.4375";
			elsif QstateRE(0) = to_sfixed(09.5000,QstateRE(0)) then
				char0RE <= "+09.5000";
			elsif QstateRE(0) = to_sfixed(09.5625,QstateRE(0)) then
				char0RE <= "+09.5625";
			elsif QstateRE(0) = to_sfixed(09.6250,QstateRE(0)) then
				char0RE <= "+09.6250";
			elsif QstateRE(0) = to_sfixed(09.6875,QstateRE(0)) then
				char0RE <= "+09.6875";
			elsif QstateRE(0) = to_sfixed(09.7500,QstateRE(0)) then
				char0RE <= "+09.7500";
			elsif QstateRE(0) = to_sfixed(09.8125,QstateRE(0)) then
				char0RE <= "+09.8125";
			elsif QstateRE(0) = to_sfixed(09.8750,QstateRE(0)) then
				char0RE <= "+09.8750";
			elsif QstateRE(0) = to_sfixed(09.9375,QstateRE(0)) then
				char0RE <= "+09.9375";
			elsif QstateRE(0) = to_sfixed(10.0000,QstateRE(0)) then
				char0RE <= "+10.0000";
			elsif QstateRE(0) = to_sfixed(10.0625,QstateRE(0)) then
				char0RE <= "+10.0625";
			elsif QstateRE(0) = to_sfixed(10.1250,QstateRE(0)) then
				char0RE <= "+10.1250";
			elsif QstateRE(0) = to_sfixed(10.1875,QstateRE(0)) then
				char0RE <= "+10.1875";
			elsif QstateRE(0) = to_sfixed(10.2500,QstateRE(0)) then
				char0RE <= "+10.2500";
			elsif QstateRE(0) = to_sfixed(10.3125,QstateRE(0)) then
				char0RE <= "+10.3125";
			elsif QstateRE(0) = to_sfixed(10.3750,QstateRE(0)) then
				char0RE <= "+10.3750";
			elsif QstateRE(0) = to_sfixed(10.4375,QstateRE(0)) then
				char0RE <= "+10.4375";
			elsif QstateRE(0) = to_sfixed(10.5000,QstateRE(0)) then
				char0RE <= "+10.5000";
			elsif QstateRE(0) = to_sfixed(10.5625,QstateRE(0)) then
				char0RE <= "+10.5625";
			elsif QstateRE(0) = to_sfixed(10.6250,QstateRE(0)) then
				char0RE <= "+10.6250";
			elsif QstateRE(0) = to_sfixed(10.6875,QstateRE(0)) then
				char0RE <= "+10.6875";
			elsif QstateRE(0) = to_sfixed(10.7500,QstateRE(0)) then
				char0RE <= "+10.7500";
			elsif QstateRE(0) = to_sfixed(10.8125,QstateRE(0)) then
				char0RE <= "+10.8125";
			elsif QstateRE(0) = to_sfixed(10.8750,QstateRE(0)) then
				char0RE <= "+10.8750";
			elsif QstateRE(0) = to_sfixed(10.9375,QstateRE(0)) then
				char0RE <= "+10.9375";
			elsif QstateRE(0) = to_sfixed(11.0000,QstateRE(0)) then
				char0RE <= "+11.0000";
			elsif QstateRE(0) = to_sfixed(11.0625,QstateRE(0)) then
				char0RE <= "+11.0625";
			elsif QstateRE(0) = to_sfixed(11.1250,QstateRE(0)) then
				char0RE <= "+11.1250";
			elsif QstateRE(0) = to_sfixed(11.1875,QstateRE(0)) then
				char0RE <= "+11.1875";
			elsif QstateRE(0) = to_sfixed(11.2500,QstateRE(0)) then
				char0RE <= "+11.2500";
			elsif QstateRE(0) = to_sfixed(11.3125,QstateRE(0)) then
				char0RE <= "+11.3125";
			elsif QstateRE(0) = to_sfixed(11.3750,QstateRE(0)) then
				char0RE <= "+11.3750";
			elsif QstateRE(0) = to_sfixed(11.4375,QstateRE(0)) then
				char0RE <= "+11.4375";
			elsif QstateRE(0) = to_sfixed(11.5000,QstateRE(0)) then
				char0RE <= "+11.5000";
			elsif QstateRE(0) = to_sfixed(11.5625,QstateRE(0)) then
				char0RE <= "+11.5625";
			elsif QstateRE(0) = to_sfixed(11.6250,QstateRE(0)) then
				char0RE <= "+11.6250";
			elsif QstateRE(0) = to_sfixed(11.6875,QstateRE(0)) then
				char0RE <= "+11.6875";
			elsif QstateRE(0) = to_sfixed(11.7500,QstateRE(0)) then
				char0RE <= "+11.7500";
			elsif QstateRE(0) = to_sfixed(11.8125,QstateRE(0)) then
				char0RE <= "+11.8125";
			elsif QstateRE(0) = to_sfixed(11.8750,QstateRE(0)) then
				char0RE <= "+11.8750";
			elsif QstateRE(0) = to_sfixed(11.9375,QstateRE(0)) then
				char0RE <= "+11.9375";
			elsif QstateRE(0) = to_sfixed(12.0000,QstateRE(0)) then
				char0RE <= "+12.0000";
			elsif QstateRE(0) = to_sfixed(12.0625,QstateRE(0)) then
				char0RE <= "+12.0625";
			elsif QstateRE(0) = to_sfixed(12.1250,QstateRE(0)) then
				char0RE <= "+12.1250";
			elsif QstateRE(0) = to_sfixed(12.1875,QstateRE(0)) then
				char0RE <= "+12.1875";
			elsif QstateRE(0) = to_sfixed(12.2500,QstateRE(0)) then
				char0RE <= "+12.2500";
			elsif QstateRE(0) = to_sfixed(12.3125,QstateRE(0)) then
				char0RE <= "+12.3125";
			elsif QstateRE(0) = to_sfixed(12.3750,QstateRE(0)) then
				char0RE <= "+12.3750";
			elsif QstateRE(0) = to_sfixed(12.4375,QstateRE(0)) then
				char0RE <= "+12.4375";
			elsif QstateRE(0) = to_sfixed(12.5000,QstateRE(0)) then
				char0RE <= "+12.5000";
			elsif QstateRE(0) = to_sfixed(12.5625,QstateRE(0)) then
				char0RE <= "+12.5625";
			elsif QstateRE(0) = to_sfixed(12.6250,QstateRE(0)) then
				char0RE <= "+12.6250";
			elsif QstateRE(0) = to_sfixed(12.6875,QstateRE(0)) then
				char0RE <= "+12.6875";
			elsif QstateRE(0) = to_sfixed(12.7500,QstateRE(0)) then
				char0RE <= "+12.7500";
			elsif QstateRE(0) = to_sfixed(12.8125,QstateRE(0)) then
				char0RE <= "+12.8125";
			elsif QstateRE(0) = to_sfixed(12.8750,QstateRE(0)) then
				char0RE <= "+12.8750";
			elsif QstateRE(0) = to_sfixed(12.9375,QstateRE(0)) then
				char0RE <= "+12.9375";
			elsif QstateRE(0) = to_sfixed(13.0000,QstateRE(0)) then
				char0RE <= "+13.0000";
			elsif QstateRE(0) = to_sfixed(13.0625,QstateRE(0)) then
				char0RE <= "+13.0625";
			elsif QstateRE(0) = to_sfixed(13.1250,QstateRE(0)) then
				char0RE <= "+13.1250";
			elsif QstateRE(0) = to_sfixed(13.1875,QstateRE(0)) then
				char0RE <= "+13.1875";
			elsif QstateRE(0) = to_sfixed(13.2500,QstateRE(0)) then
				char0RE <= "+13.2500";
			elsif QstateRE(0) = to_sfixed(13.3125,QstateRE(0)) then
				char0RE <= "+13.3125";
			elsif QstateRE(0) = to_sfixed(13.3750,QstateRE(0)) then
				char0RE <= "+13.3750";
			elsif QstateRE(0) = to_sfixed(13.4375,QstateRE(0)) then
				char0RE <= "+13.4375";
			elsif QstateRE(0) = to_sfixed(13.5000,QstateRE(0)) then
				char0RE <= "+13.5000";
			elsif QstateRE(0) = to_sfixed(13.5625,QstateRE(0)) then
				char0RE <= "+13.5625";
			elsif QstateRE(0) = to_sfixed(13.6250,QstateRE(0)) then
				char0RE <= "+13.6250";
			elsif QstateRE(0) = to_sfixed(13.6875,QstateRE(0)) then
				char0RE <= "+13.6875";
			elsif QstateRE(0) = to_sfixed(13.7500,QstateRE(0)) then
				char0RE <= "+13.7500";
			elsif QstateRE(0) = to_sfixed(13.8125,QstateRE(0)) then
				char0RE <= "+13.8125";
			elsif QstateRE(0) = to_sfixed(13.8750,QstateRE(0)) then
				char0RE <= "+13.8750";
			elsif QstateRE(0) = to_sfixed(13.9375,QstateRE(0)) then
				char0RE <= "+13.9375";
			elsif QstateRE(0) = to_sfixed(14.0000,QstateRE(0)) then
				char0RE <= "+14.0000";
			elsif QstateRE(0) = to_sfixed(14.0625,QstateRE(0)) then
				char0RE <= "+14.0625";
			elsif QstateRE(0) = to_sfixed(14.1250,QstateRE(0)) then
				char0RE <= "+14.1250";
			elsif QstateRE(0) = to_sfixed(14.1875,QstateRE(0)) then
				char0RE <= "+14.1875";
			elsif QstateRE(0) = to_sfixed(14.2500,QstateRE(0)) then
				char0RE <= "+14.2500";
			elsif QstateRE(0) = to_sfixed(14.3125,QstateRE(0)) then
				char0RE <= "+14.3125";
			elsif QstateRE(0) = to_sfixed(14.3750,QstateRE(0)) then
				char0RE <= "+14.3750";
			elsif QstateRE(0) = to_sfixed(14.4375,QstateRE(0)) then
				char0RE <= "+14.4375";
			elsif QstateRE(0) = to_sfixed(14.5000,QstateRE(0)) then
				char0RE <= "+14.5000";
			elsif QstateRE(0) = to_sfixed(14.5625,QstateRE(0)) then
				char0RE <= "+14.5625";
			elsif QstateRE(0) = to_sfixed(14.6250,QstateRE(0)) then
				char0RE <= "+14.6250";
			elsif QstateRE(0) = to_sfixed(14.6875,QstateRE(0)) then
				char0RE <= "+14.6875";
			elsif QstateRE(0) = to_sfixed(14.7500,QstateRE(0)) then
				char0RE <= "+14.7500";
			elsif QstateRE(0) = to_sfixed(14.8125,QstateRE(0)) then
				char0RE <= "+14.8125";
			elsif QstateRE(0) = to_sfixed(14.8750,QstateRE(0)) then
				char0RE <= "+14.8750";
			elsif QstateRE(0) = to_sfixed(14.9375,QstateRE(0)) then
				char0RE <= "+14.9375";
			elsif QstateRE(0) = to_sfixed(15.0000,QstateRE(0)) then
				char0RE <= "+15.0000";
			elsif QstateRE(0) = to_sfixed(15.0625,QstateRE(0)) then
				char0RE <= "+15.0625";
			elsif QstateRE(0) = to_sfixed(15.1250,QstateRE(0)) then
				char0RE <= "+15.1250";
			elsif QstateRE(0) = to_sfixed(15.1875,QstateRE(0)) then
				char0RE <= "+15.1875";
			elsif QstateRE(0) = to_sfixed(15.2500,QstateRE(0)) then
				char0RE <= "+15.2500";
			elsif QstateRE(0) = to_sfixed(15.3125,QstateRE(0)) then
				char0RE <= "+15.3125";
			elsif QstateRE(0) = to_sfixed(15.3750,QstateRE(0)) then
				char0RE <= "+15.3750";
			elsif QstateRE(0) = to_sfixed(15.4375,QstateRE(0)) then
				char0RE <= "+15.4375";
			elsif QstateRE(0) = to_sfixed(15.5000,QstateRE(0)) then
				char0RE <= "+15.5000";
			elsif QstateRE(0) = to_sfixed(15.5625,QstateRE(0)) then
				char0RE <= "+15.5625";
			elsif QstateRE(0) = to_sfixed(15.6250,QstateRE(0)) then
				char0RE <= "+15.6250";
			elsif QstateRE(0) = to_sfixed(15.6875,QstateRE(0)) then
				char0RE <= "+15.6875";
			elsif QstateRE(0) = to_sfixed(15.7500,QstateRE(0)) then
				char0RE <= "+15.7500";
			elsif QstateRE(0) = to_sfixed(15.8125,QstateRE(0)) then
				char0RE <= "+15.8125";
			elsif QstateRE(0) = to_sfixed(15.8750,QstateRE(0)) then
				char0RE <= "+15.8750";
			elsif QstateRE(0) = to_sfixed(15.9375,QstateRE(0)) then
				char0RE <= "+15.9375";
			end if;
			if QstateIM(0) = to_sfixed(-15.9375,QstateIM(0)) then
				char0IM <= "-15.9375";
			elsif QstateIM(0) = to_sfixed(-15.8750,QstateIM(0)) then
				char0IM <= "-15.8750";
			elsif QstateIM(0) = to_sfixed(-15.8125,QstateIM(0)) then
				char0IM <= "-15.8125";
			elsif QstateIM(0) = to_sfixed(-15.7500,QstateIM(0)) then
				char0IM <= "-15.7500";
			elsif QstateIM(0) = to_sfixed(-15.6875,QstateIM(0)) then
				char0IM <= "-15.6875";
			elsif QstateIM(0) = to_sfixed(-15.6250,QstateIM(0)) then
				char0IM <= "-15.6250";
			elsif QstateIM(0) = to_sfixed(-15.5625,QstateIM(0)) then
				char0IM <= "-15.5625";
			elsif QstateIM(0) = to_sfixed(-15.5000,QstateIM(0)) then
				char0IM <= "-15.5000";
			elsif QstateIM(0) = to_sfixed(-15.4375,QstateIM(0)) then
				char0IM <= "-15.4375";
			elsif QstateIM(0) = to_sfixed(-15.3750,QstateIM(0)) then
				char0IM <= "-15.3750";
			elsif QstateIM(0) = to_sfixed(-15.3125,QstateIM(0)) then
				char0IM <= "-15.3125";
			elsif QstateIM(0) = to_sfixed(-15.2500,QstateIM(0)) then
				char0IM <= "-15.2500";
			elsif QstateIM(0) = to_sfixed(-15.1875,QstateIM(0)) then
				char0IM <= "-15.1875";
			elsif QstateIM(0) = to_sfixed(-15.1250,QstateIM(0)) then
				char0IM <= "-15.1250";
			elsif QstateIM(0) = to_sfixed(-15.0625,QstateIM(0)) then
				char0IM <= "-15.0625";
			elsif QstateIM(0) = to_sfixed(-15.0000,QstateIM(0)) then
				char0IM <= "-15.0000";
			elsif QstateIM(0) = to_sfixed(-14.9375,QstateIM(0)) then
				char0IM <= "-14.9375";
			elsif QstateIM(0) = to_sfixed(-14.8750,QstateIM(0)) then
				char0IM <= "-14.8750";
			elsif QstateIM(0) = to_sfixed(-14.8125,QstateIM(0)) then
				char0IM <= "-14.8125";
			elsif QstateIM(0) = to_sfixed(-14.7500,QstateIM(0)) then
				char0IM <= "-14.7500";
			elsif QstateIM(0) = to_sfixed(-14.6875,QstateIM(0)) then
				char0IM <= "-14.6875";
			elsif QstateIM(0) = to_sfixed(-14.6250,QstateIM(0)) then
				char0IM <= "-14.6250";
			elsif QstateIM(0) = to_sfixed(-14.5625,QstateIM(0)) then
				char0IM <= "-14.5625";
			elsif QstateIM(0) = to_sfixed(-14.5000,QstateIM(0)) then
				char0IM <= "-14.5000";
			elsif QstateIM(0) = to_sfixed(-14.4375,QstateIM(0)) then
				char0IM <= "-14.4375";
			elsif QstateIM(0) = to_sfixed(-14.3750,QstateIM(0)) then
				char0IM <= "-14.3750";
			elsif QstateIM(0) = to_sfixed(-14.3125,QstateIM(0)) then
				char0IM <= "-14.3125";
			elsif QstateIM(0) = to_sfixed(-14.2500,QstateIM(0)) then
				char0IM <= "-14.2500";
			elsif QstateIM(0) = to_sfixed(-14.1875,QstateIM(0)) then
				char0IM <= "-14.1875";
			elsif QstateIM(0) = to_sfixed(-14.1250,QstateIM(0)) then
				char0IM <= "-14.1250";
			elsif QstateIM(0) = to_sfixed(-14.0625,QstateIM(0)) then
				char0IM <= "-14.0625";
			elsif QstateIM(0) = to_sfixed(-14.0000,QstateIM(0)) then
				char0IM <= "-14.0000";
			elsif QstateIM(0) = to_sfixed(-13.9375,QstateIM(0)) then
				char0IM <= "-13.9375";
			elsif QstateIM(0) = to_sfixed(-13.8750,QstateIM(0)) then
				char0IM <= "-13.8750";
			elsif QstateIM(0) = to_sfixed(-13.8125,QstateIM(0)) then
				char0IM <= "-13.8125";
			elsif QstateIM(0) = to_sfixed(-13.7500,QstateIM(0)) then
				char0IM <= "-13.7500";
			elsif QstateIM(0) = to_sfixed(-13.6875,QstateIM(0)) then
				char0IM <= "-13.6875";
			elsif QstateIM(0) = to_sfixed(-13.6250,QstateIM(0)) then
				char0IM <= "-13.6250";
			elsif QstateIM(0) = to_sfixed(-13.5625,QstateIM(0)) then
				char0IM <= "-13.5625";
			elsif QstateIM(0) = to_sfixed(-13.5000,QstateIM(0)) then
				char0IM <= "-13.5000";
			elsif QstateIM(0) = to_sfixed(-13.4375,QstateIM(0)) then
				char0IM <= "-13.4375";
			elsif QstateIM(0) = to_sfixed(-13.3750,QstateIM(0)) then
				char0IM <= "-13.3750";
			elsif QstateIM(0) = to_sfixed(-13.3125,QstateIM(0)) then
				char0IM <= "-13.3125";
			elsif QstateIM(0) = to_sfixed(-13.2500,QstateIM(0)) then
				char0IM <= "-13.2500";
			elsif QstateIM(0) = to_sfixed(-13.1875,QstateIM(0)) then
				char0IM <= "-13.1875";
			elsif QstateIM(0) = to_sfixed(-13.1250,QstateIM(0)) then
				char0IM <= "-13.1250";
			elsif QstateIM(0) = to_sfixed(-13.0625,QstateIM(0)) then
				char0IM <= "-13.0625";
			elsif QstateIM(0) = to_sfixed(-13.0000,QstateIM(0)) then
				char0IM <= "-13.0000";
			elsif QstateIM(0) = to_sfixed(-12.9375,QstateIM(0)) then
				char0IM <= "-12.9375";
			elsif QstateIM(0) = to_sfixed(-12.8750,QstateIM(0)) then
				char0IM <= "-12.8750";
			elsif QstateIM(0) = to_sfixed(-12.8125,QstateIM(0)) then
				char0IM <= "-12.8125";
			elsif QstateIM(0) = to_sfixed(-12.7500,QstateIM(0)) then
				char0IM <= "-12.7500";
			elsif QstateIM(0) = to_sfixed(-12.6875,QstateIM(0)) then
				char0IM <= "-12.6875";
			elsif QstateIM(0) = to_sfixed(-12.6250,QstateIM(0)) then
				char0IM <= "-12.6250";
			elsif QstateIM(0) = to_sfixed(-12.5625,QstateIM(0)) then
				char0IM <= "-12.5625";
			elsif QstateIM(0) = to_sfixed(-12.5000,QstateIM(0)) then
				char0IM <= "-12.5000";
			elsif QstateIM(0) = to_sfixed(-12.4375,QstateIM(0)) then
				char0IM <= "-12.4375";
			elsif QstateIM(0) = to_sfixed(-12.3750,QstateIM(0)) then
				char0IM <= "-12.3750";
			elsif QstateIM(0) = to_sfixed(-12.3125,QstateIM(0)) then
				char0IM <= "-12.3125";
			elsif QstateIM(0) = to_sfixed(-12.2500,QstateIM(0)) then
				char0IM <= "-12.2500";
			elsif QstateIM(0) = to_sfixed(-12.1875,QstateIM(0)) then
				char0IM <= "-12.1875";
			elsif QstateIM(0) = to_sfixed(-12.1250,QstateIM(0)) then
				char0IM <= "-12.1250";
			elsif QstateIM(0) = to_sfixed(-12.0625,QstateIM(0)) then
				char0IM <= "-12.0625";
			elsif QstateIM(0) = to_sfixed(-12.0000,QstateIM(0)) then
				char0IM <= "-12.0000";
			elsif QstateIM(0) = to_sfixed(-11.9375,QstateIM(0)) then
				char0IM <= "-11.9375";
			elsif QstateIM(0) = to_sfixed(-11.8750,QstateIM(0)) then
				char0IM <= "-11.8750";
			elsif QstateIM(0) = to_sfixed(-11.8125,QstateIM(0)) then
				char0IM <= "-11.8125";
			elsif QstateIM(0) = to_sfixed(-11.7500,QstateIM(0)) then
				char0IM <= "-11.7500";
			elsif QstateIM(0) = to_sfixed(-11.6875,QstateIM(0)) then
				char0IM <= "-11.6875";
			elsif QstateIM(0) = to_sfixed(-11.6250,QstateIM(0)) then
				char0IM <= "-11.6250";
			elsif QstateIM(0) = to_sfixed(-11.5625,QstateIM(0)) then
				char0IM <= "-11.5625";
			elsif QstateIM(0) = to_sfixed(-11.5000,QstateIM(0)) then
				char0IM <= "-11.5000";
			elsif QstateIM(0) = to_sfixed(-11.4375,QstateIM(0)) then
				char0IM <= "-11.4375";
			elsif QstateIM(0) = to_sfixed(-11.3750,QstateIM(0)) then
				char0IM <= "-11.3750";
			elsif QstateIM(0) = to_sfixed(-11.3125,QstateIM(0)) then
				char0IM <= "-11.3125";
			elsif QstateIM(0) = to_sfixed(-11.2500,QstateIM(0)) then
				char0IM <= "-11.2500";
			elsif QstateIM(0) = to_sfixed(-11.1875,QstateIM(0)) then
				char0IM <= "-11.1875";
			elsif QstateIM(0) = to_sfixed(-11.1250,QstateIM(0)) then
				char0IM <= "-11.1250";
			elsif QstateIM(0) = to_sfixed(-11.0625,QstateIM(0)) then
				char0IM <= "-11.0625";
			elsif QstateIM(0) = to_sfixed(-11.0000,QstateIM(0)) then
				char0IM <= "-11.0000";
			elsif QstateIM(0) = to_sfixed(-10.9375,QstateIM(0)) then
				char0IM <= "-10.9375";
			elsif QstateIM(0) = to_sfixed(-10.8750,QstateIM(0)) then
				char0IM <= "-10.8750";
			elsif QstateIM(0) = to_sfixed(-10.8125,QstateIM(0)) then
				char0IM <= "-10.8125";
			elsif QstateIM(0) = to_sfixed(-10.7500,QstateIM(0)) then
				char0IM <= "-10.7500";
			elsif QstateIM(0) = to_sfixed(-10.6875,QstateIM(0)) then
				char0IM <= "-10.6875";
			elsif QstateIM(0) = to_sfixed(-10.6250,QstateIM(0)) then
				char0IM <= "-10.6250";
			elsif QstateIM(0) = to_sfixed(-10.5625,QstateIM(0)) then
				char0IM <= "-10.5625";
			elsif QstateIM(0) = to_sfixed(-10.5000,QstateIM(0)) then
				char0IM <= "-10.5000";
			elsif QstateIM(0) = to_sfixed(-10.4375,QstateIM(0)) then
				char0IM <= "-10.4375";
			elsif QstateIM(0) = to_sfixed(-10.3750,QstateIM(0)) then
				char0IM <= "-10.3750";
			elsif QstateIM(0) = to_sfixed(-10.3125,QstateIM(0)) then
				char0IM <= "-10.3125";
			elsif QstateIM(0) = to_sfixed(-10.2500,QstateIM(0)) then
				char0IM <= "-10.2500";
			elsif QstateIM(0) = to_sfixed(-10.1875,QstateIM(0)) then
				char0IM <= "-10.1875";
			elsif QstateIM(0) = to_sfixed(-10.1250,QstateIM(0)) then
				char0IM <= "-10.1250";
			elsif QstateIM(0) = to_sfixed(-10.0625,QstateIM(0)) then
				char0IM <= "-10.0625";
			elsif QstateIM(0) = to_sfixed(-10.0000,QstateIM(0)) then
				char0IM <= "-10.0000";
			elsif QstateIM(0) = to_sfixed(-9.9375,QstateIM(0)) then
				char0IM <= "--9.9375";
			elsif QstateIM(0) = to_sfixed(-9.8750,QstateIM(0)) then
				char0IM <= "--9.8750";
			elsif QstateIM(0) = to_sfixed(-9.8125,QstateIM(0)) then
				char0IM <= "--9.8125";
			elsif QstateIM(0) = to_sfixed(-9.7500,QstateIM(0)) then
				char0IM <= "--9.7500";
			elsif QstateIM(0) = to_sfixed(-9.6875,QstateIM(0)) then
				char0IM <= "--9.6875";
			elsif QstateIM(0) = to_sfixed(-9.6250,QstateIM(0)) then
				char0IM <= "--9.6250";
			elsif QstateIM(0) = to_sfixed(-9.5625,QstateIM(0)) then
				char0IM <= "--9.5625";
			elsif QstateIM(0) = to_sfixed(-9.5000,QstateIM(0)) then
				char0IM <= "--9.5000";
			elsif QstateIM(0) = to_sfixed(-9.4375,QstateIM(0)) then
				char0IM <= "--9.4375";
			elsif QstateIM(0) = to_sfixed(-9.3750,QstateIM(0)) then
				char0IM <= "--9.3750";
			elsif QstateIM(0) = to_sfixed(-9.3125,QstateIM(0)) then
				char0IM <= "--9.3125";
			elsif QstateIM(0) = to_sfixed(-9.2500,QstateIM(0)) then
				char0IM <= "--9.2500";
			elsif QstateIM(0) = to_sfixed(-9.1875,QstateIM(0)) then
				char0IM <= "--9.1875";
			elsif QstateIM(0) = to_sfixed(-9.1250,QstateIM(0)) then
				char0IM <= "--9.1250";
			elsif QstateIM(0) = to_sfixed(-9.0625,QstateIM(0)) then
				char0IM <= "--9.0625";
			elsif QstateIM(0) = to_sfixed(-9.0000,QstateIM(0)) then
				char0IM <= "--9.0000";
			elsif QstateIM(0) = to_sfixed(-8.9375,QstateIM(0)) then
				char0IM <= "--8.9375";
			elsif QstateIM(0) = to_sfixed(-8.8750,QstateIM(0)) then
				char0IM <= "--8.8750";
			elsif QstateIM(0) = to_sfixed(-8.8125,QstateIM(0)) then
				char0IM <= "--8.8125";
			elsif QstateIM(0) = to_sfixed(-8.7500,QstateIM(0)) then
				char0IM <= "--8.7500";
			elsif QstateIM(0) = to_sfixed(-8.6875,QstateIM(0)) then
				char0IM <= "--8.6875";
			elsif QstateIM(0) = to_sfixed(-8.6250,QstateIM(0)) then
				char0IM <= "--8.6250";
			elsif QstateIM(0) = to_sfixed(-8.5625,QstateIM(0)) then
				char0IM <= "--8.5625";
			elsif QstateIM(0) = to_sfixed(-8.5000,QstateIM(0)) then
				char0IM <= "--8.5000";
			elsif QstateIM(0) = to_sfixed(-8.4375,QstateIM(0)) then
				char0IM <= "--8.4375";
			elsif QstateIM(0) = to_sfixed(-8.3750,QstateIM(0)) then
				char0IM <= "--8.3750";
			elsif QstateIM(0) = to_sfixed(-8.3125,QstateIM(0)) then
				char0IM <= "--8.3125";
			elsif QstateIM(0) = to_sfixed(-8.2500,QstateIM(0)) then
				char0IM <= "--8.2500";
			elsif QstateIM(0) = to_sfixed(-8.1875,QstateIM(0)) then
				char0IM <= "--8.1875";
			elsif QstateIM(0) = to_sfixed(-8.1250,QstateIM(0)) then
				char0IM <= "--8.1250";
			elsif QstateIM(0) = to_sfixed(-8.0625,QstateIM(0)) then
				char0IM <= "--8.0625";
			elsif QstateIM(0) = to_sfixed(-8.0000,QstateIM(0)) then
				char0IM <= "--8.0000";
			elsif QstateIM(0) = to_sfixed(-7.9375,QstateIM(0)) then
				char0IM <= "--7.9375";
			elsif QstateIM(0) = to_sfixed(-7.8750,QstateIM(0)) then
				char0IM <= "--7.8750";
			elsif QstateIM(0) = to_sfixed(-7.8125,QstateIM(0)) then
				char0IM <= "--7.8125";
			elsif QstateIM(0) = to_sfixed(-7.7500,QstateIM(0)) then
				char0IM <= "--7.7500";
			elsif QstateIM(0) = to_sfixed(-7.6875,QstateIM(0)) then
				char0IM <= "--7.6875";
			elsif QstateIM(0) = to_sfixed(-7.6250,QstateIM(0)) then
				char0IM <= "--7.6250";
			elsif QstateIM(0) = to_sfixed(-7.5625,QstateIM(0)) then
				char0IM <= "--7.5625";
			elsif QstateIM(0) = to_sfixed(-7.5000,QstateIM(0)) then
				char0IM <= "--7.5000";
			elsif QstateIM(0) = to_sfixed(-7.4375,QstateIM(0)) then
				char0IM <= "--7.4375";
			elsif QstateIM(0) = to_sfixed(-7.3750,QstateIM(0)) then
				char0IM <= "--7.3750";
			elsif QstateIM(0) = to_sfixed(-7.3125,QstateIM(0)) then
				char0IM <= "--7.3125";
			elsif QstateIM(0) = to_sfixed(-7.2500,QstateIM(0)) then
				char0IM <= "--7.2500";
			elsif QstateIM(0) = to_sfixed(-7.1875,QstateIM(0)) then
				char0IM <= "--7.1875";
			elsif QstateIM(0) = to_sfixed(-7.1250,QstateIM(0)) then
				char0IM <= "--7.1250";
			elsif QstateIM(0) = to_sfixed(-7.0625,QstateIM(0)) then
				char0IM <= "--7.0625";
			elsif QstateIM(0) = to_sfixed(-7.0000,QstateIM(0)) then
				char0IM <= "--7.0000";
			elsif QstateIM(0) = to_sfixed(-6.9375,QstateIM(0)) then
				char0IM <= "--6.9375";
			elsif QstateIM(0) = to_sfixed(-6.8750,QstateIM(0)) then
				char0IM <= "--6.8750";
			elsif QstateIM(0) = to_sfixed(-6.8125,QstateIM(0)) then
				char0IM <= "--6.8125";
			elsif QstateIM(0) = to_sfixed(-6.7500,QstateIM(0)) then
				char0IM <= "--6.7500";
			elsif QstateIM(0) = to_sfixed(-6.6875,QstateIM(0)) then
				char0IM <= "--6.6875";
			elsif QstateIM(0) = to_sfixed(-6.6250,QstateIM(0)) then
				char0IM <= "--6.6250";
			elsif QstateIM(0) = to_sfixed(-6.5625,QstateIM(0)) then
				char0IM <= "--6.5625";
			elsif QstateIM(0) = to_sfixed(-6.5000,QstateIM(0)) then
				char0IM <= "--6.5000";
			elsif QstateIM(0) = to_sfixed(-6.4375,QstateIM(0)) then
				char0IM <= "--6.4375";
			elsif QstateIM(0) = to_sfixed(-6.3750,QstateIM(0)) then
				char0IM <= "--6.3750";
			elsif QstateIM(0) = to_sfixed(-6.3125,QstateIM(0)) then
				char0IM <= "--6.3125";
			elsif QstateIM(0) = to_sfixed(-6.2500,QstateIM(0)) then
				char0IM <= "--6.2500";
			elsif QstateIM(0) = to_sfixed(-6.1875,QstateIM(0)) then
				char0IM <= "--6.1875";
			elsif QstateIM(0) = to_sfixed(-6.1250,QstateIM(0)) then
				char0IM <= "--6.1250";
			elsif QstateIM(0) = to_sfixed(-6.0625,QstateIM(0)) then
				char0IM <= "--6.0625";
			elsif QstateIM(0) = to_sfixed(-6.0000,QstateIM(0)) then
				char0IM <= "--6.0000";
			elsif QstateIM(0) = to_sfixed(-5.9375,QstateIM(0)) then
				char0IM <= "--5.9375";
			elsif QstateIM(0) = to_sfixed(-5.8750,QstateIM(0)) then
				char0IM <= "--5.8750";
			elsif QstateIM(0) = to_sfixed(-5.8125,QstateIM(0)) then
				char0IM <= "--5.8125";
			elsif QstateIM(0) = to_sfixed(-5.7500,QstateIM(0)) then
				char0IM <= "--5.7500";
			elsif QstateIM(0) = to_sfixed(-5.6875,QstateIM(0)) then
				char0IM <= "--5.6875";
			elsif QstateIM(0) = to_sfixed(-5.6250,QstateIM(0)) then
				char0IM <= "--5.6250";
			elsif QstateIM(0) = to_sfixed(-5.5625,QstateIM(0)) then
				char0IM <= "--5.5625";
			elsif QstateIM(0) = to_sfixed(-5.5000,QstateIM(0)) then
				char0IM <= "--5.5000";
			elsif QstateIM(0) = to_sfixed(-5.4375,QstateIM(0)) then
				char0IM <= "--5.4375";
			elsif QstateIM(0) = to_sfixed(-5.3750,QstateIM(0)) then
				char0IM <= "--5.3750";
			elsif QstateIM(0) = to_sfixed(-5.3125,QstateIM(0)) then
				char0IM <= "--5.3125";
			elsif QstateIM(0) = to_sfixed(-5.2500,QstateIM(0)) then
				char0IM <= "--5.2500";
			elsif QstateIM(0) = to_sfixed(-5.1875,QstateIM(0)) then
				char0IM <= "--5.1875";
			elsif QstateIM(0) = to_sfixed(-5.1250,QstateIM(0)) then
				char0IM <= "--5.1250";
			elsif QstateIM(0) = to_sfixed(-5.0625,QstateIM(0)) then
				char0IM <= "--5.0625";
			elsif QstateIM(0) = to_sfixed(-5.0000,QstateIM(0)) then
				char0IM <= "--5.0000";
			elsif QstateIM(0) = to_sfixed(-4.9375,QstateIM(0)) then
				char0IM <= "--4.9375";
			elsif QstateIM(0) = to_sfixed(-4.8750,QstateIM(0)) then
				char0IM <= "--4.8750";
			elsif QstateIM(0) = to_sfixed(-4.8125,QstateIM(0)) then
				char0IM <= "--4.8125";
			elsif QstateIM(0) = to_sfixed(-4.7500,QstateIM(0)) then
				char0IM <= "--4.7500";
			elsif QstateIM(0) = to_sfixed(-4.6875,QstateIM(0)) then
				char0IM <= "--4.6875";
			elsif QstateIM(0) = to_sfixed(-4.6250,QstateIM(0)) then
				char0IM <= "--4.6250";
			elsif QstateIM(0) = to_sfixed(-4.5625,QstateIM(0)) then
				char0IM <= "--4.5625";
			elsif QstateIM(0) = to_sfixed(-4.5000,QstateIM(0)) then
				char0IM <= "--4.5000";
			elsif QstateIM(0) = to_sfixed(-4.4375,QstateIM(0)) then
				char0IM <= "--4.4375";
			elsif QstateIM(0) = to_sfixed(-4.3750,QstateIM(0)) then
				char0IM <= "--4.3750";
			elsif QstateIM(0) = to_sfixed(-4.3125,QstateIM(0)) then
				char0IM <= "--4.3125";
			elsif QstateIM(0) = to_sfixed(-4.2500,QstateIM(0)) then
				char0IM <= "--4.2500";
			elsif QstateIM(0) = to_sfixed(-4.1875,QstateIM(0)) then
				char0IM <= "--4.1875";
			elsif QstateIM(0) = to_sfixed(-4.1250,QstateIM(0)) then
				char0IM <= "--4.1250";
			elsif QstateIM(0) = to_sfixed(-4.0625,QstateIM(0)) then
				char0IM <= "--4.0625";
			elsif QstateIM(0) = to_sfixed(-4.0000,QstateIM(0)) then
				char0IM <= "--4.0000";
			elsif QstateIM(0) = to_sfixed(-3.9375,QstateIM(0)) then
				char0IM <= "--3.9375";
			elsif QstateIM(0) = to_sfixed(-3.8750,QstateIM(0)) then
				char0IM <= "--3.8750";
			elsif QstateIM(0) = to_sfixed(-3.8125,QstateIM(0)) then
				char0IM <= "--3.8125";
			elsif QstateIM(0) = to_sfixed(-3.7500,QstateIM(0)) then
				char0IM <= "--3.7500";
			elsif QstateIM(0) = to_sfixed(-3.6875,QstateIM(0)) then
				char0IM <= "--3.6875";
			elsif QstateIM(0) = to_sfixed(-3.6250,QstateIM(0)) then
				char0IM <= "--3.6250";
			elsif QstateIM(0) = to_sfixed(-3.5625,QstateIM(0)) then
				char0IM <= "--3.5625";
			elsif QstateIM(0) = to_sfixed(-3.5000,QstateIM(0)) then
				char0IM <= "--3.5000";
			elsif QstateIM(0) = to_sfixed(-3.4375,QstateIM(0)) then
				char0IM <= "--3.4375";
			elsif QstateIM(0) = to_sfixed(-3.3750,QstateIM(0)) then
				char0IM <= "--3.3750";
			elsif QstateIM(0) = to_sfixed(-3.3125,QstateIM(0)) then
				char0IM <= "--3.3125";
			elsif QstateIM(0) = to_sfixed(-3.2500,QstateIM(0)) then
				char0IM <= "--3.2500";
			elsif QstateIM(0) = to_sfixed(-3.1875,QstateIM(0)) then
				char0IM <= "--3.1875";
			elsif QstateIM(0) = to_sfixed(-3.1250,QstateIM(0)) then
				char0IM <= "--3.1250";
			elsif QstateIM(0) = to_sfixed(-3.0625,QstateIM(0)) then
				char0IM <= "--3.0625";
			elsif QstateIM(0) = to_sfixed(-3.0000,QstateIM(0)) then
				char0IM <= "--3.0000";
			elsif QstateIM(0) = to_sfixed(-2.9375,QstateIM(0)) then
				char0IM <= "--2.9375";
			elsif QstateIM(0) = to_sfixed(-2.8750,QstateIM(0)) then
				char0IM <= "--2.8750";
			elsif QstateIM(0) = to_sfixed(-2.8125,QstateIM(0)) then
				char0IM <= "--2.8125";
			elsif QstateIM(0) = to_sfixed(-2.7500,QstateIM(0)) then
				char0IM <= "--2.7500";
			elsif QstateIM(0) = to_sfixed(-2.6875,QstateIM(0)) then
				char0IM <= "--2.6875";
			elsif QstateIM(0) = to_sfixed(-2.6250,QstateIM(0)) then
				char0IM <= "--2.6250";
			elsif QstateIM(0) = to_sfixed(-2.5625,QstateIM(0)) then
				char0IM <= "--2.5625";
			elsif QstateIM(0) = to_sfixed(-2.5000,QstateIM(0)) then
				char0IM <= "--2.5000";
			elsif QstateIM(0) = to_sfixed(-2.4375,QstateIM(0)) then
				char0IM <= "--2.4375";
			elsif QstateIM(0) = to_sfixed(-2.3750,QstateIM(0)) then
				char0IM <= "--2.3750";
			elsif QstateIM(0) = to_sfixed(-2.3125,QstateIM(0)) then
				char0IM <= "--2.3125";
			elsif QstateIM(0) = to_sfixed(-2.2500,QstateIM(0)) then
				char0IM <= "--2.2500";
			elsif QstateIM(0) = to_sfixed(-2.1875,QstateIM(0)) then
				char0IM <= "--2.1875";
			elsif QstateIM(0) = to_sfixed(-2.1250,QstateIM(0)) then
				char0IM <= "--2.1250";
			elsif QstateIM(0) = to_sfixed(-2.0625,QstateIM(0)) then
				char0IM <= "--2.0625";
			elsif QstateIM(0) = to_sfixed(-2.0000,QstateIM(0)) then
				char0IM <= "--2.0000";
			elsif QstateIM(0) = to_sfixed(-1.9375,QstateIM(0)) then
				char0IM <= "--1.9375";
			elsif QstateIM(0) = to_sfixed(-1.8750,QstateIM(0)) then
				char0IM <= "--1.8750";
			elsif QstateIM(0) = to_sfixed(-1.8125,QstateIM(0)) then
				char0IM <= "--1.8125";
			elsif QstateIM(0) = to_sfixed(-1.7500,QstateIM(0)) then
				char0IM <= "--1.7500";
			elsif QstateIM(0) = to_sfixed(-1.6875,QstateIM(0)) then
				char0IM <= "--1.6875";
			elsif QstateIM(0) = to_sfixed(-1.6250,QstateIM(0)) then
				char0IM <= "--1.6250";
			elsif QstateIM(0) = to_sfixed(-1.5625,QstateIM(0)) then
				char0IM <= "--1.5625";
			elsif QstateIM(0) = to_sfixed(-1.5000,QstateIM(0)) then
				char0IM <= "--1.5000";
			elsif QstateIM(0) = to_sfixed(-1.4375,QstateIM(0)) then
				char0IM <= "--1.4375";
			elsif QstateIM(0) = to_sfixed(-1.3750,QstateIM(0)) then
				char0IM <= "--1.3750";
			elsif QstateIM(0) = to_sfixed(-1.3125,QstateIM(0)) then
				char0IM <= "--1.3125";
			elsif QstateIM(0) = to_sfixed(-1.2500,QstateIM(0)) then
				char0IM <= "--1.2500";
			elsif QstateIM(0) = to_sfixed(-1.1875,QstateIM(0)) then
				char0IM <= "--1.1875";
			elsif QstateIM(0) = to_sfixed(-1.1250,QstateIM(0)) then
				char0IM <= "--1.1250";
			elsif QstateIM(0) = to_sfixed(-1.0625,QstateIM(0)) then
				char0IM <= "--1.0625";
			elsif QstateIM(0) = to_sfixed(-1.0000,QstateIM(0)) then
				char0IM <= "--1.0000";
			elsif QstateIM(0) = to_sfixed(-0.9375,QstateIM(0)) then
				char0IM <= "--0.9375";
			elsif QstateIM(0) = to_sfixed(-0.8750,QstateIM(0)) then
				char0IM <= "--0.8750";
			elsif QstateIM(0) = to_sfixed(-0.8125,QstateIM(0)) then
				char0IM <= "--0.8125";
			elsif QstateIM(0) = to_sfixed(-0.7500,QstateIM(0)) then
				char0IM <= "--0.7500";
			elsif QstateIM(0) = to_sfixed(-0.6875,QstateIM(0)) then
				char0IM <= "--0.6875";
			elsif QstateIM(0) = to_sfixed(-0.6250,QstateIM(0)) then
				char0IM <= "--0.6250";
			elsif QstateIM(0) = to_sfixed(-0.5625,QstateIM(0)) then
				char0IM <= "--0.5625";
			elsif QstateIM(0) = to_sfixed(-0.5000,QstateIM(0)) then
				char0IM <= "--0.5000";
			elsif QstateIM(0) = to_sfixed(-0.4375,QstateIM(0)) then
				char0IM <= "--0.4375";
			elsif QstateIM(0) = to_sfixed(-0.3750,QstateIM(0)) then
				char0IM <= "--0.3750";
			elsif QstateIM(0) = to_sfixed(-0.3125,QstateIM(0)) then
				char0IM <= "--0.3125";
			elsif QstateIM(0) = to_sfixed(-0.2500,QstateIM(0)) then
				char0IM <= "--0.2500";
			elsif QstateIM(0) = to_sfixed(-0.1875,QstateIM(0)) then
				char0IM <= "--0.1875";
			elsif QstateIM(0) = to_sfixed(-0.1250,QstateIM(0)) then
				char0IM <= "--0.1250";
			elsif QstateIM(0) = to_sfixed(-0.0625,QstateIM(0)) then
				char0IM <= "--0.0625";
			elsif QstateIM(0) = to_sfixed(00.0000,QstateIM(0)) then
				char0IM <= "+00.0000";
			elsif QstateIM(0) = to_sfixed(00.0625,QstateIM(0)) then
				char0IM <= "+00.0625";
			elsif QstateIM(0) = to_sfixed(00.1250,QstateIM(0)) then
				char0IM <= "+00.1250";
			elsif QstateIM(0) = to_sfixed(00.1875,QstateIM(0)) then
				char0IM <= "+00.1875";
			elsif QstateIM(0) = to_sfixed(00.2500,QstateIM(0)) then
				char0IM <= "+00.2500";
			elsif QstateIM(0) = to_sfixed(00.3125,QstateIM(0)) then
				char0IM <= "+00.3125";
			elsif QstateIM(0) = to_sfixed(00.3750,QstateIM(0)) then
				char0IM <= "+00.3750";
			elsif QstateIM(0) = to_sfixed(00.4375,QstateIM(0)) then
				char0IM <= "+00.4375";
			elsif QstateIM(0) = to_sfixed(00.5000,QstateIM(0)) then
				char0IM <= "+00.5000";
			elsif QstateIM(0) = to_sfixed(00.5625,QstateIM(0)) then
				char0IM <= "+00.5625";
			elsif QstateIM(0) = to_sfixed(00.6250,QstateIM(0)) then
				char0IM <= "+00.6250";
			elsif QstateIM(0) = to_sfixed(00.6875,QstateIM(0)) then
				char0IM <= "+00.6875";
			elsif QstateIM(0) = to_sfixed(00.7500,QstateIM(0)) then
				char0IM <= "+00.7500";
			elsif QstateIM(0) = to_sfixed(00.8125,QstateIM(0)) then
				char0IM <= "+00.8125";
			elsif QstateIM(0) = to_sfixed(00.8750,QstateIM(0)) then
				char0IM <= "+00.8750";
			elsif QstateIM(0) = to_sfixed(00.9375,QstateIM(0)) then
				char0IM <= "+00.9375";
			elsif QstateIM(0) = to_sfixed(01.0000,QstateIM(0)) then
				char0IM <= "+01.0000";
			elsif QstateIM(0) = to_sfixed(01.0625,QstateIM(0)) then
				char0IM <= "+01.0625";
			elsif QstateIM(0) = to_sfixed(01.1250,QstateIM(0)) then
				char0IM <= "+01.1250";
			elsif QstateIM(0) = to_sfixed(01.1875,QstateIM(0)) then
				char0IM <= "+01.1875";
			elsif QstateIM(0) = to_sfixed(01.2500,QstateIM(0)) then
				char0IM <= "+01.2500";
			elsif QstateIM(0) = to_sfixed(01.3125,QstateIM(0)) then
				char0IM <= "+01.3125";
			elsif QstateIM(0) = to_sfixed(01.3750,QstateIM(0)) then
				char0IM <= "+01.3750";
			elsif QstateIM(0) = to_sfixed(01.4375,QstateIM(0)) then
				char0IM <= "+01.4375";
			elsif QstateIM(0) = to_sfixed(01.5000,QstateIM(0)) then
				char0IM <= "+01.5000";
			elsif QstateIM(0) = to_sfixed(01.5625,QstateIM(0)) then
				char0IM <= "+01.5625";
			elsif QstateIM(0) = to_sfixed(01.6250,QstateIM(0)) then
				char0IM <= "+01.6250";
			elsif QstateIM(0) = to_sfixed(01.6875,QstateIM(0)) then
				char0IM <= "+01.6875";
			elsif QstateIM(0) = to_sfixed(01.7500,QstateIM(0)) then
				char0IM <= "+01.7500";
			elsif QstateIM(0) = to_sfixed(01.8125,QstateIM(0)) then
				char0IM <= "+01.8125";
			elsif QstateIM(0) = to_sfixed(01.8750,QstateIM(0)) then
				char0IM <= "+01.8750";
			elsif QstateIM(0) = to_sfixed(01.9375,QstateIM(0)) then
				char0IM <= "+01.9375";
			elsif QstateIM(0) = to_sfixed(02.0000,QstateIM(0)) then
				char0IM <= "+02.0000";
			elsif QstateIM(0) = to_sfixed(02.0625,QstateIM(0)) then
				char0IM <= "+02.0625";
			elsif QstateIM(0) = to_sfixed(02.1250,QstateIM(0)) then
				char0IM <= "+02.1250";
			elsif QstateIM(0) = to_sfixed(02.1875,QstateIM(0)) then
				char0IM <= "+02.1875";
			elsif QstateIM(0) = to_sfixed(02.2500,QstateIM(0)) then
				char0IM <= "+02.2500";
			elsif QstateIM(0) = to_sfixed(02.3125,QstateIM(0)) then
				char0IM <= "+02.3125";
			elsif QstateIM(0) = to_sfixed(02.3750,QstateIM(0)) then
				char0IM <= "+02.3750";
			elsif QstateIM(0) = to_sfixed(02.4375,QstateIM(0)) then
				char0IM <= "+02.4375";
			elsif QstateIM(0) = to_sfixed(02.5000,QstateIM(0)) then
				char0IM <= "+02.5000";
			elsif QstateIM(0) = to_sfixed(02.5625,QstateIM(0)) then
				char0IM <= "+02.5625";
			elsif QstateIM(0) = to_sfixed(02.6250,QstateIM(0)) then
				char0IM <= "+02.6250";
			elsif QstateIM(0) = to_sfixed(02.6875,QstateIM(0)) then
				char0IM <= "+02.6875";
			elsif QstateIM(0) = to_sfixed(02.7500,QstateIM(0)) then
				char0IM <= "+02.7500";
			elsif QstateIM(0) = to_sfixed(02.8125,QstateIM(0)) then
				char0IM <= "+02.8125";
			elsif QstateIM(0) = to_sfixed(02.8750,QstateIM(0)) then
				char0IM <= "+02.8750";
			elsif QstateIM(0) = to_sfixed(02.9375,QstateIM(0)) then
				char0IM <= "+02.9375";
			elsif QstateIM(0) = to_sfixed(03.0000,QstateIM(0)) then
				char0IM <= "+03.0000";
			elsif QstateIM(0) = to_sfixed(03.0625,QstateIM(0)) then
				char0IM <= "+03.0625";
			elsif QstateIM(0) = to_sfixed(03.1250,QstateIM(0)) then
				char0IM <= "+03.1250";
			elsif QstateIM(0) = to_sfixed(03.1875,QstateIM(0)) then
				char0IM <= "+03.1875";
			elsif QstateIM(0) = to_sfixed(03.2500,QstateIM(0)) then
				char0IM <= "+03.2500";
			elsif QstateIM(0) = to_sfixed(03.3125,QstateIM(0)) then
				char0IM <= "+03.3125";
			elsif QstateIM(0) = to_sfixed(03.3750,QstateIM(0)) then
				char0IM <= "+03.3750";
			elsif QstateIM(0) = to_sfixed(03.4375,QstateIM(0)) then
				char0IM <= "+03.4375";
			elsif QstateIM(0) = to_sfixed(03.5000,QstateIM(0)) then
				char0IM <= "+03.5000";
			elsif QstateIM(0) = to_sfixed(03.5625,QstateIM(0)) then
				char0IM <= "+03.5625";
			elsif QstateIM(0) = to_sfixed(03.6250,QstateIM(0)) then
				char0IM <= "+03.6250";
			elsif QstateIM(0) = to_sfixed(03.6875,QstateIM(0)) then
				char0IM <= "+03.6875";
			elsif QstateIM(0) = to_sfixed(03.7500,QstateIM(0)) then
				char0IM <= "+03.7500";
			elsif QstateIM(0) = to_sfixed(03.8125,QstateIM(0)) then
				char0IM <= "+03.8125";
			elsif QstateIM(0) = to_sfixed(03.8750,QstateIM(0)) then
				char0IM <= "+03.8750";
			elsif QstateIM(0) = to_sfixed(03.9375,QstateIM(0)) then
				char0IM <= "+03.9375";
			elsif QstateIM(0) = to_sfixed(04.0000,QstateIM(0)) then
				char0IM <= "+04.0000";
			elsif QstateIM(0) = to_sfixed(04.0625,QstateIM(0)) then
				char0IM <= "+04.0625";
			elsif QstateIM(0) = to_sfixed(04.1250,QstateIM(0)) then
				char0IM <= "+04.1250";
			elsif QstateIM(0) = to_sfixed(04.1875,QstateIM(0)) then
				char0IM <= "+04.1875";
			elsif QstateIM(0) = to_sfixed(04.2500,QstateIM(0)) then
				char0IM <= "+04.2500";
			elsif QstateIM(0) = to_sfixed(04.3125,QstateIM(0)) then
				char0IM <= "+04.3125";
			elsif QstateIM(0) = to_sfixed(04.3750,QstateIM(0)) then
				char0IM <= "+04.3750";
			elsif QstateIM(0) = to_sfixed(04.4375,QstateIM(0)) then
				char0IM <= "+04.4375";
			elsif QstateIM(0) = to_sfixed(04.5000,QstateIM(0)) then
				char0IM <= "+04.5000";
			elsif QstateIM(0) = to_sfixed(04.5625,QstateIM(0)) then
				char0IM <= "+04.5625";
			elsif QstateIM(0) = to_sfixed(04.6250,QstateIM(0)) then
				char0IM <= "+04.6250";
			elsif QstateIM(0) = to_sfixed(04.6875,QstateIM(0)) then
				char0IM <= "+04.6875";
			elsif QstateIM(0) = to_sfixed(04.7500,QstateIM(0)) then
				char0IM <= "+04.7500";
			elsif QstateIM(0) = to_sfixed(04.8125,QstateIM(0)) then
				char0IM <= "+04.8125";
			elsif QstateIM(0) = to_sfixed(04.8750,QstateIM(0)) then
				char0IM <= "+04.8750";
			elsif QstateIM(0) = to_sfixed(04.9375,QstateIM(0)) then
				char0IM <= "+04.9375";
			elsif QstateIM(0) = to_sfixed(05.0000,QstateIM(0)) then
				char0IM <= "+05.0000";
			elsif QstateIM(0) = to_sfixed(05.0625,QstateIM(0)) then
				char0IM <= "+05.0625";
			elsif QstateIM(0) = to_sfixed(05.1250,QstateIM(0)) then
				char0IM <= "+05.1250";
			elsif QstateIM(0) = to_sfixed(05.1875,QstateIM(0)) then
				char0IM <= "+05.1875";
			elsif QstateIM(0) = to_sfixed(05.2500,QstateIM(0)) then
				char0IM <= "+05.2500";
			elsif QstateIM(0) = to_sfixed(05.3125,QstateIM(0)) then
				char0IM <= "+05.3125";
			elsif QstateIM(0) = to_sfixed(05.3750,QstateIM(0)) then
				char0IM <= "+05.3750";
			elsif QstateIM(0) = to_sfixed(05.4375,QstateIM(0)) then
				char0IM <= "+05.4375";
			elsif QstateIM(0) = to_sfixed(05.5000,QstateIM(0)) then
				char0IM <= "+05.5000";
			elsif QstateIM(0) = to_sfixed(05.5625,QstateIM(0)) then
				char0IM <= "+05.5625";
			elsif QstateIM(0) = to_sfixed(05.6250,QstateIM(0)) then
				char0IM <= "+05.6250";
			elsif QstateIM(0) = to_sfixed(05.6875,QstateIM(0)) then
				char0IM <= "+05.6875";
			elsif QstateIM(0) = to_sfixed(05.7500,QstateIM(0)) then
				char0IM <= "+05.7500";
			elsif QstateIM(0) = to_sfixed(05.8125,QstateIM(0)) then
				char0IM <= "+05.8125";
			elsif QstateIM(0) = to_sfixed(05.8750,QstateIM(0)) then
				char0IM <= "+05.8750";
			elsif QstateIM(0) = to_sfixed(05.9375,QstateIM(0)) then
				char0IM <= "+05.9375";
			elsif QstateIM(0) = to_sfixed(06.0000,QstateIM(0)) then
				char0IM <= "+06.0000";
			elsif QstateIM(0) = to_sfixed(06.0625,QstateIM(0)) then
				char0IM <= "+06.0625";
			elsif QstateIM(0) = to_sfixed(06.1250,QstateIM(0)) then
				char0IM <= "+06.1250";
			elsif QstateIM(0) = to_sfixed(06.1875,QstateIM(0)) then
				char0IM <= "+06.1875";
			elsif QstateIM(0) = to_sfixed(06.2500,QstateIM(0)) then
				char0IM <= "+06.2500";
			elsif QstateIM(0) = to_sfixed(06.3125,QstateIM(0)) then
				char0IM <= "+06.3125";
			elsif QstateIM(0) = to_sfixed(06.3750,QstateIM(0)) then
				char0IM <= "+06.3750";
			elsif QstateIM(0) = to_sfixed(06.4375,QstateIM(0)) then
				char0IM <= "+06.4375";
			elsif QstateIM(0) = to_sfixed(06.5000,QstateIM(0)) then
				char0IM <= "+06.5000";
			elsif QstateIM(0) = to_sfixed(06.5625,QstateIM(0)) then
				char0IM <= "+06.5625";
			elsif QstateIM(0) = to_sfixed(06.6250,QstateIM(0)) then
				char0IM <= "+06.6250";
			elsif QstateIM(0) = to_sfixed(06.6875,QstateIM(0)) then
				char0IM <= "+06.6875";
			elsif QstateIM(0) = to_sfixed(06.7500,QstateIM(0)) then
				char0IM <= "+06.7500";
			elsif QstateIM(0) = to_sfixed(06.8125,QstateIM(0)) then
				char0IM <= "+06.8125";
			elsif QstateIM(0) = to_sfixed(06.8750,QstateIM(0)) then
				char0IM <= "+06.8750";
			elsif QstateIM(0) = to_sfixed(06.9375,QstateIM(0)) then
				char0IM <= "+06.9375";
			elsif QstateIM(0) = to_sfixed(07.0000,QstateIM(0)) then
				char0IM <= "+07.0000";
			elsif QstateIM(0) = to_sfixed(07.0625,QstateIM(0)) then
				char0IM <= "+07.0625";
			elsif QstateIM(0) = to_sfixed(07.1250,QstateIM(0)) then
				char0IM <= "+07.1250";
			elsif QstateIM(0) = to_sfixed(07.1875,QstateIM(0)) then
				char0IM <= "+07.1875";
			elsif QstateIM(0) = to_sfixed(07.2500,QstateIM(0)) then
				char0IM <= "+07.2500";
			elsif QstateIM(0) = to_sfixed(07.3125,QstateIM(0)) then
				char0IM <= "+07.3125";
			elsif QstateIM(0) = to_sfixed(07.3750,QstateIM(0)) then
				char0IM <= "+07.3750";
			elsif QstateIM(0) = to_sfixed(07.4375,QstateIM(0)) then
				char0IM <= "+07.4375";
			elsif QstateIM(0) = to_sfixed(07.5000,QstateIM(0)) then
				char0IM <= "+07.5000";
			elsif QstateIM(0) = to_sfixed(07.5625,QstateIM(0)) then
				char0IM <= "+07.5625";
			elsif QstateIM(0) = to_sfixed(07.6250,QstateIM(0)) then
				char0IM <= "+07.6250";
			elsif QstateIM(0) = to_sfixed(07.6875,QstateIM(0)) then
				char0IM <= "+07.6875";
			elsif QstateIM(0) = to_sfixed(07.7500,QstateIM(0)) then
				char0IM <= "+07.7500";
			elsif QstateIM(0) = to_sfixed(07.8125,QstateIM(0)) then
				char0IM <= "+07.8125";
			elsif QstateIM(0) = to_sfixed(07.8750,QstateIM(0)) then
				char0IM <= "+07.8750";
			elsif QstateIM(0) = to_sfixed(07.9375,QstateIM(0)) then
				char0IM <= "+07.9375";
			elsif QstateIM(0) = to_sfixed(08.0000,QstateIM(0)) then
				char0IM <= "+08.0000";
			elsif QstateIM(0) = to_sfixed(08.0625,QstateIM(0)) then
				char0IM <= "+08.0625";
			elsif QstateIM(0) = to_sfixed(08.1250,QstateIM(0)) then
				char0IM <= "+08.1250";
			elsif QstateIM(0) = to_sfixed(08.1875,QstateIM(0)) then
				char0IM <= "+08.1875";
			elsif QstateIM(0) = to_sfixed(08.2500,QstateIM(0)) then
				char0IM <= "+08.2500";
			elsif QstateIM(0) = to_sfixed(08.3125,QstateIM(0)) then
				char0IM <= "+08.3125";
			elsif QstateIM(0) = to_sfixed(08.3750,QstateIM(0)) then
				char0IM <= "+08.3750";
			elsif QstateIM(0) = to_sfixed(08.4375,QstateIM(0)) then
				char0IM <= "+08.4375";
			elsif QstateIM(0) = to_sfixed(08.5000,QstateIM(0)) then
				char0IM <= "+08.5000";
			elsif QstateIM(0) = to_sfixed(08.5625,QstateIM(0)) then
				char0IM <= "+08.5625";
			elsif QstateIM(0) = to_sfixed(08.6250,QstateIM(0)) then
				char0IM <= "+08.6250";
			elsif QstateIM(0) = to_sfixed(08.6875,QstateIM(0)) then
				char0IM <= "+08.6875";
			elsif QstateIM(0) = to_sfixed(08.7500,QstateIM(0)) then
				char0IM <= "+08.7500";
			elsif QstateIM(0) = to_sfixed(08.8125,QstateIM(0)) then
				char0IM <= "+08.8125";
			elsif QstateIM(0) = to_sfixed(08.8750,QstateIM(0)) then
				char0IM <= "+08.8750";
			elsif QstateIM(0) = to_sfixed(08.9375,QstateIM(0)) then
				char0IM <= "+08.9375";
			elsif QstateIM(0) = to_sfixed(09.0000,QstateIM(0)) then
				char0IM <= "+09.0000";
			elsif QstateIM(0) = to_sfixed(09.0625,QstateIM(0)) then
				char0IM <= "+09.0625";
			elsif QstateIM(0) = to_sfixed(09.1250,QstateIM(0)) then
				char0IM <= "+09.1250";
			elsif QstateIM(0) = to_sfixed(09.1875,QstateIM(0)) then
				char0IM <= "+09.1875";
			elsif QstateIM(0) = to_sfixed(09.2500,QstateIM(0)) then
				char0IM <= "+09.2500";
			elsif QstateIM(0) = to_sfixed(09.3125,QstateIM(0)) then
				char0IM <= "+09.3125";
			elsif QstateIM(0) = to_sfixed(09.3750,QstateIM(0)) then
				char0IM <= "+09.3750";
			elsif QstateIM(0) = to_sfixed(09.4375,QstateIM(0)) then
				char0IM <= "+09.4375";
			elsif QstateIM(0) = to_sfixed(09.5000,QstateIM(0)) then
				char0IM <= "+09.5000";
			elsif QstateIM(0) = to_sfixed(09.5625,QstateIM(0)) then
				char0IM <= "+09.5625";
			elsif QstateIM(0) = to_sfixed(09.6250,QstateIM(0)) then
				char0IM <= "+09.6250";
			elsif QstateIM(0) = to_sfixed(09.6875,QstateIM(0)) then
				char0IM <= "+09.6875";
			elsif QstateIM(0) = to_sfixed(09.7500,QstateIM(0)) then
				char0IM <= "+09.7500";
			elsif QstateIM(0) = to_sfixed(09.8125,QstateIM(0)) then
				char0IM <= "+09.8125";
			elsif QstateIM(0) = to_sfixed(09.8750,QstateIM(0)) then
				char0IM <= "+09.8750";
			elsif QstateIM(0) = to_sfixed(09.9375,QstateIM(0)) then
				char0IM <= "+09.9375";
			elsif QstateIM(0) = to_sfixed(10.0000,QstateIM(0)) then
				char0IM <= "+10.0000";
			elsif QstateIM(0) = to_sfixed(10.0625,QstateIM(0)) then
				char0IM <= "+10.0625";
			elsif QstateIM(0) = to_sfixed(10.1250,QstateIM(0)) then
				char0IM <= "+10.1250";
			elsif QstateIM(0) = to_sfixed(10.1875,QstateIM(0)) then
				char0IM <= "+10.1875";
			elsif QstateIM(0) = to_sfixed(10.2500,QstateIM(0)) then
				char0IM <= "+10.2500";
			elsif QstateIM(0) = to_sfixed(10.3125,QstateIM(0)) then
				char0IM <= "+10.3125";
			elsif QstateIM(0) = to_sfixed(10.3750,QstateIM(0)) then
				char0IM <= "+10.3750";
			elsif QstateIM(0) = to_sfixed(10.4375,QstateIM(0)) then
				char0IM <= "+10.4375";
			elsif QstateIM(0) = to_sfixed(10.5000,QstateIM(0)) then
				char0IM <= "+10.5000";
			elsif QstateIM(0) = to_sfixed(10.5625,QstateIM(0)) then
				char0IM <= "+10.5625";
			elsif QstateIM(0) = to_sfixed(10.6250,QstateIM(0)) then
				char0IM <= "+10.6250";
			elsif QstateIM(0) = to_sfixed(10.6875,QstateIM(0)) then
				char0IM <= "+10.6875";
			elsif QstateIM(0) = to_sfixed(10.7500,QstateIM(0)) then
				char0IM <= "+10.7500";
			elsif QstateIM(0) = to_sfixed(10.8125,QstateIM(0)) then
				char0IM <= "+10.8125";
			elsif QstateIM(0) = to_sfixed(10.8750,QstateIM(0)) then
				char0IM <= "+10.8750";
			elsif QstateIM(0) = to_sfixed(10.9375,QstateIM(0)) then
				char0IM <= "+10.9375";
			elsif QstateIM(0) = to_sfixed(11.0000,QstateIM(0)) then
				char0IM <= "+11.0000";
			elsif QstateIM(0) = to_sfixed(11.0625,QstateIM(0)) then
				char0IM <= "+11.0625";
			elsif QstateIM(0) = to_sfixed(11.1250,QstateIM(0)) then
				char0IM <= "+11.1250";
			elsif QstateIM(0) = to_sfixed(11.1875,QstateIM(0)) then
				char0IM <= "+11.1875";
			elsif QstateIM(0) = to_sfixed(11.2500,QstateIM(0)) then
				char0IM <= "+11.2500";
			elsif QstateIM(0) = to_sfixed(11.3125,QstateIM(0)) then
				char0IM <= "+11.3125";
			elsif QstateIM(0) = to_sfixed(11.3750,QstateIM(0)) then
				char0IM <= "+11.3750";
			elsif QstateIM(0) = to_sfixed(11.4375,QstateIM(0)) then
				char0IM <= "+11.4375";
			elsif QstateIM(0) = to_sfixed(11.5000,QstateIM(0)) then
				char0IM <= "+11.5000";
			elsif QstateIM(0) = to_sfixed(11.5625,QstateIM(0)) then
				char0IM <= "+11.5625";
			elsif QstateIM(0) = to_sfixed(11.6250,QstateIM(0)) then
				char0IM <= "+11.6250";
			elsif QstateIM(0) = to_sfixed(11.6875,QstateIM(0)) then
				char0IM <= "+11.6875";
			elsif QstateIM(0) = to_sfixed(11.7500,QstateIM(0)) then
				char0IM <= "+11.7500";
			elsif QstateIM(0) = to_sfixed(11.8125,QstateIM(0)) then
				char0IM <= "+11.8125";
			elsif QstateIM(0) = to_sfixed(11.8750,QstateIM(0)) then
				char0IM <= "+11.8750";
			elsif QstateIM(0) = to_sfixed(11.9375,QstateIM(0)) then
				char0IM <= "+11.9375";
			elsif QstateIM(0) = to_sfixed(12.0000,QstateIM(0)) then
				char0IM <= "+12.0000";
			elsif QstateIM(0) = to_sfixed(12.0625,QstateIM(0)) then
				char0IM <= "+12.0625";
			elsif QstateIM(0) = to_sfixed(12.1250,QstateIM(0)) then
				char0IM <= "+12.1250";
			elsif QstateIM(0) = to_sfixed(12.1875,QstateIM(0)) then
				char0IM <= "+12.1875";
			elsif QstateIM(0) = to_sfixed(12.2500,QstateIM(0)) then
				char0IM <= "+12.2500";
			elsif QstateIM(0) = to_sfixed(12.3125,QstateIM(0)) then
				char0IM <= "+12.3125";
			elsif QstateIM(0) = to_sfixed(12.3750,QstateIM(0)) then
				char0IM <= "+12.3750";
			elsif QstateIM(0) = to_sfixed(12.4375,QstateIM(0)) then
				char0IM <= "+12.4375";
			elsif QstateIM(0) = to_sfixed(12.5000,QstateIM(0)) then
				char0IM <= "+12.5000";
			elsif QstateIM(0) = to_sfixed(12.5625,QstateIM(0)) then
				char0IM <= "+12.5625";
			elsif QstateIM(0) = to_sfixed(12.6250,QstateIM(0)) then
				char0IM <= "+12.6250";
			elsif QstateIM(0) = to_sfixed(12.6875,QstateIM(0)) then
				char0IM <= "+12.6875";
			elsif QstateIM(0) = to_sfixed(12.7500,QstateIM(0)) then
				char0IM <= "+12.7500";
			elsif QstateIM(0) = to_sfixed(12.8125,QstateIM(0)) then
				char0IM <= "+12.8125";
			elsif QstateIM(0) = to_sfixed(12.8750,QstateIM(0)) then
				char0IM <= "+12.8750";
			elsif QstateIM(0) = to_sfixed(12.9375,QstateIM(0)) then
				char0IM <= "+12.9375";
			elsif QstateIM(0) = to_sfixed(13.0000,QstateIM(0)) then
				char0IM <= "+13.0000";
			elsif QstateIM(0) = to_sfixed(13.0625,QstateIM(0)) then
				char0IM <= "+13.0625";
			elsif QstateIM(0) = to_sfixed(13.1250,QstateIM(0)) then
				char0IM <= "+13.1250";
			elsif QstateIM(0) = to_sfixed(13.1875,QstateIM(0)) then
				char0IM <= "+13.1875";
			elsif QstateIM(0) = to_sfixed(13.2500,QstateIM(0)) then
				char0IM <= "+13.2500";
			elsif QstateIM(0) = to_sfixed(13.3125,QstateIM(0)) then
				char0IM <= "+13.3125";
			elsif QstateIM(0) = to_sfixed(13.3750,QstateIM(0)) then
				char0IM <= "+13.3750";
			elsif QstateIM(0) = to_sfixed(13.4375,QstateIM(0)) then
				char0IM <= "+13.4375";
			elsif QstateIM(0) = to_sfixed(13.5000,QstateIM(0)) then
				char0IM <= "+13.5000";
			elsif QstateIM(0) = to_sfixed(13.5625,QstateIM(0)) then
				char0IM <= "+13.5625";
			elsif QstateIM(0) = to_sfixed(13.6250,QstateIM(0)) then
				char0IM <= "+13.6250";
			elsif QstateIM(0) = to_sfixed(13.6875,QstateIM(0)) then
				char0IM <= "+13.6875";
			elsif QstateIM(0) = to_sfixed(13.7500,QstateIM(0)) then
				char0IM <= "+13.7500";
			elsif QstateIM(0) = to_sfixed(13.8125,QstateIM(0)) then
				char0IM <= "+13.8125";
			elsif QstateIM(0) = to_sfixed(13.8750,QstateIM(0)) then
				char0IM <= "+13.8750";
			elsif QstateIM(0) = to_sfixed(13.9375,QstateIM(0)) then
				char0IM <= "+13.9375";
			elsif QstateIM(0) = to_sfixed(14.0000,QstateIM(0)) then
				char0IM <= "+14.0000";
			elsif QstateIM(0) = to_sfixed(14.0625,QstateIM(0)) then
				char0IM <= "+14.0625";
			elsif QstateIM(0) = to_sfixed(14.1250,QstateIM(0)) then
				char0IM <= "+14.1250";
			elsif QstateIM(0) = to_sfixed(14.1875,QstateIM(0)) then
				char0IM <= "+14.1875";
			elsif QstateIM(0) = to_sfixed(14.2500,QstateIM(0)) then
				char0IM <= "+14.2500";
			elsif QstateIM(0) = to_sfixed(14.3125,QstateIM(0)) then
				char0IM <= "+14.3125";
			elsif QstateIM(0) = to_sfixed(14.3750,QstateIM(0)) then
				char0IM <= "+14.3750";
			elsif QstateIM(0) = to_sfixed(14.4375,QstateIM(0)) then
				char0IM <= "+14.4375";
			elsif QstateIM(0) = to_sfixed(14.5000,QstateIM(0)) then
				char0IM <= "+14.5000";
			elsif QstateIM(0) = to_sfixed(14.5625,QstateIM(0)) then
				char0IM <= "+14.5625";
			elsif QstateIM(0) = to_sfixed(14.6250,QstateIM(0)) then
				char0IM <= "+14.6250";
			elsif QstateIM(0) = to_sfixed(14.6875,QstateIM(0)) then
				char0IM <= "+14.6875";
			elsif QstateIM(0) = to_sfixed(14.7500,QstateIM(0)) then
				char0IM <= "+14.7500";
			elsif QstateIM(0) = to_sfixed(14.8125,QstateIM(0)) then
				char0IM <= "+14.8125";
			elsif QstateIM(0) = to_sfixed(14.8750,QstateIM(0)) then
				char0IM <= "+14.8750";
			elsif QstateIM(0) = to_sfixed(14.9375,QstateIM(0)) then
				char0IM <= "+14.9375";
			elsif QstateIM(0) = to_sfixed(15.0000,QstateIM(0)) then
				char0IM <= "+15.0000";
			elsif QstateIM(0) = to_sfixed(15.0625,QstateIM(0)) then
				char0IM <= "+15.0625";
			elsif QstateIM(0) = to_sfixed(15.1250,QstateIM(0)) then
				char0IM <= "+15.1250";
			elsif QstateIM(0) = to_sfixed(15.1875,QstateIM(0)) then
				char0IM <= "+15.1875";
			elsif QstateIM(0) = to_sfixed(15.2500,QstateIM(0)) then
				char0IM <= "+15.2500";
			elsif QstateIM(0) = to_sfixed(15.3125,QstateIM(0)) then
				char0IM <= "+15.3125";
			elsif QstateIM(0) = to_sfixed(15.3750,QstateIM(0)) then
				char0IM <= "+15.3750";
			elsif QstateIM(0) = to_sfixed(15.4375,QstateIM(0)) then
				char0IM <= "+15.4375";
			elsif QstateIM(0) = to_sfixed(15.5000,QstateIM(0)) then
				char0IM <= "+15.5000";
			elsif QstateIM(0) = to_sfixed(15.5625,QstateIM(0)) then
				char0IM <= "+15.5625";
			elsif QstateIM(0) = to_sfixed(15.6250,QstateIM(0)) then
				char0IM <= "+15.6250";
			elsif QstateIM(0) = to_sfixed(15.6875,QstateIM(0)) then
				char0IM <= "+15.6875";
			elsif QstateIM(0) = to_sfixed(15.7500,QstateIM(0)) then
				char0IM <= "+15.7500";
			elsif QstateIM(0) = to_sfixed(15.8125,QstateIM(0)) then
				char0IM <= "+15.8125";
			elsif QstateIM(0) = to_sfixed(15.8750,QstateIM(0)) then
				char0IM <= "+15.8750";
			elsif QstateIM(0) = to_sfixed(15.9375,QstateIM(0)) then
				char0IM <= "+15.9375";
			end if;
			if QstateRE(1) = to_sfixed(-15.9375,QstateRE(1)) then
				char1RE <= "-15.9375";
			elsif QstateRE(1) = to_sfixed(-15.8750,QstateRE(1)) then
				char1RE <= "-15.8750";
			elsif QstateRE(1) = to_sfixed(-15.8125,QstateRE(1)) then
				char1RE <= "-15.8125";
			elsif QstateRE(1) = to_sfixed(-15.7500,QstateRE(1)) then
				char1RE <= "-15.7500";
			elsif QstateRE(1) = to_sfixed(-15.6875,QstateRE(1)) then
				char1RE <= "-15.6875";
			elsif QstateRE(1) = to_sfixed(-15.6250,QstateRE(1)) then
				char1RE <= "-15.6250";
			elsif QstateRE(1) = to_sfixed(-15.5625,QstateRE(1)) then
				char1RE <= "-15.5625";
			elsif QstateRE(1) = to_sfixed(-15.5000,QstateRE(1)) then
				char1RE <= "-15.5000";
			elsif QstateRE(1) = to_sfixed(-15.4375,QstateRE(1)) then
				char1RE <= "-15.4375";
			elsif QstateRE(1) = to_sfixed(-15.3750,QstateRE(1)) then
				char1RE <= "-15.3750";
			elsif QstateRE(1) = to_sfixed(-15.3125,QstateRE(1)) then
				char1RE <= "-15.3125";
			elsif QstateRE(1) = to_sfixed(-15.2500,QstateRE(1)) then
				char1RE <= "-15.2500";
			elsif QstateRE(1) = to_sfixed(-15.1875,QstateRE(1)) then
				char1RE <= "-15.1875";
			elsif QstateRE(1) = to_sfixed(-15.1250,QstateRE(1)) then
				char1RE <= "-15.1250";
			elsif QstateRE(1) = to_sfixed(-15.0625,QstateRE(1)) then
				char1RE <= "-15.0625";
			elsif QstateRE(1) = to_sfixed(-15.0000,QstateRE(1)) then
				char1RE <= "-15.0000";
			elsif QstateRE(1) = to_sfixed(-14.9375,QstateRE(1)) then
				char1RE <= "-14.9375";
			elsif QstateRE(1) = to_sfixed(-14.8750,QstateRE(1)) then
				char1RE <= "-14.8750";
			elsif QstateRE(1) = to_sfixed(-14.8125,QstateRE(1)) then
				char1RE <= "-14.8125";
			elsif QstateRE(1) = to_sfixed(-14.7500,QstateRE(1)) then
				char1RE <= "-14.7500";
			elsif QstateRE(1) = to_sfixed(-14.6875,QstateRE(1)) then
				char1RE <= "-14.6875";
			elsif QstateRE(1) = to_sfixed(-14.6250,QstateRE(1)) then
				char1RE <= "-14.6250";
			elsif QstateRE(1) = to_sfixed(-14.5625,QstateRE(1)) then
				char1RE <= "-14.5625";
			elsif QstateRE(1) = to_sfixed(-14.5000,QstateRE(1)) then
				char1RE <= "-14.5000";
			elsif QstateRE(1) = to_sfixed(-14.4375,QstateRE(1)) then
				char1RE <= "-14.4375";
			elsif QstateRE(1) = to_sfixed(-14.3750,QstateRE(1)) then
				char1RE <= "-14.3750";
			elsif QstateRE(1) = to_sfixed(-14.3125,QstateRE(1)) then
				char1RE <= "-14.3125";
			elsif QstateRE(1) = to_sfixed(-14.2500,QstateRE(1)) then
				char1RE <= "-14.2500";
			elsif QstateRE(1) = to_sfixed(-14.1875,QstateRE(1)) then
				char1RE <= "-14.1875";
			elsif QstateRE(1) = to_sfixed(-14.1250,QstateRE(1)) then
				char1RE <= "-14.1250";
			elsif QstateRE(1) = to_sfixed(-14.0625,QstateRE(1)) then
				char1RE <= "-14.0625";
			elsif QstateRE(1) = to_sfixed(-14.0000,QstateRE(1)) then
				char1RE <= "-14.0000";
			elsif QstateRE(1) = to_sfixed(-13.9375,QstateRE(1)) then
				char1RE <= "-13.9375";
			elsif QstateRE(1) = to_sfixed(-13.8750,QstateRE(1)) then
				char1RE <= "-13.8750";
			elsif QstateRE(1) = to_sfixed(-13.8125,QstateRE(1)) then
				char1RE <= "-13.8125";
			elsif QstateRE(1) = to_sfixed(-13.7500,QstateRE(1)) then
				char1RE <= "-13.7500";
			elsif QstateRE(1) = to_sfixed(-13.6875,QstateRE(1)) then
				char1RE <= "-13.6875";
			elsif QstateRE(1) = to_sfixed(-13.6250,QstateRE(1)) then
				char1RE <= "-13.6250";
			elsif QstateRE(1) = to_sfixed(-13.5625,QstateRE(1)) then
				char1RE <= "-13.5625";
			elsif QstateRE(1) = to_sfixed(-13.5000,QstateRE(1)) then
				char1RE <= "-13.5000";
			elsif QstateRE(1) = to_sfixed(-13.4375,QstateRE(1)) then
				char1RE <= "-13.4375";
			elsif QstateRE(1) = to_sfixed(-13.3750,QstateRE(1)) then
				char1RE <= "-13.3750";
			elsif QstateRE(1) = to_sfixed(-13.3125,QstateRE(1)) then
				char1RE <= "-13.3125";
			elsif QstateRE(1) = to_sfixed(-13.2500,QstateRE(1)) then
				char1RE <= "-13.2500";
			elsif QstateRE(1) = to_sfixed(-13.1875,QstateRE(1)) then
				char1RE <= "-13.1875";
			elsif QstateRE(1) = to_sfixed(-13.1250,QstateRE(1)) then
				char1RE <= "-13.1250";
			elsif QstateRE(1) = to_sfixed(-13.0625,QstateRE(1)) then
				char1RE <= "-13.0625";
			elsif QstateRE(1) = to_sfixed(-13.0000,QstateRE(1)) then
				char1RE <= "-13.0000";
			elsif QstateRE(1) = to_sfixed(-12.9375,QstateRE(1)) then
				char1RE <= "-12.9375";
			elsif QstateRE(1) = to_sfixed(-12.8750,QstateRE(1)) then
				char1RE <= "-12.8750";
			elsif QstateRE(1) = to_sfixed(-12.8125,QstateRE(1)) then
				char1RE <= "-12.8125";
			elsif QstateRE(1) = to_sfixed(-12.7500,QstateRE(1)) then
				char1RE <= "-12.7500";
			elsif QstateRE(1) = to_sfixed(-12.6875,QstateRE(1)) then
				char1RE <= "-12.6875";
			elsif QstateRE(1) = to_sfixed(-12.6250,QstateRE(1)) then
				char1RE <= "-12.6250";
			elsif QstateRE(1) = to_sfixed(-12.5625,QstateRE(1)) then
				char1RE <= "-12.5625";
			elsif QstateRE(1) = to_sfixed(-12.5000,QstateRE(1)) then
				char1RE <= "-12.5000";
			elsif QstateRE(1) = to_sfixed(-12.4375,QstateRE(1)) then
				char1RE <= "-12.4375";
			elsif QstateRE(1) = to_sfixed(-12.3750,QstateRE(1)) then
				char1RE <= "-12.3750";
			elsif QstateRE(1) = to_sfixed(-12.3125,QstateRE(1)) then
				char1RE <= "-12.3125";
			elsif QstateRE(1) = to_sfixed(-12.2500,QstateRE(1)) then
				char1RE <= "-12.2500";
			elsif QstateRE(1) = to_sfixed(-12.1875,QstateRE(1)) then
				char1RE <= "-12.1875";
			elsif QstateRE(1) = to_sfixed(-12.1250,QstateRE(1)) then
				char1RE <= "-12.1250";
			elsif QstateRE(1) = to_sfixed(-12.0625,QstateRE(1)) then
				char1RE <= "-12.0625";
			elsif QstateRE(1) = to_sfixed(-12.0000,QstateRE(1)) then
				char1RE <= "-12.0000";
			elsif QstateRE(1) = to_sfixed(-11.9375,QstateRE(1)) then
				char1RE <= "-11.9375";
			elsif QstateRE(1) = to_sfixed(-11.8750,QstateRE(1)) then
				char1RE <= "-11.8750";
			elsif QstateRE(1) = to_sfixed(-11.8125,QstateRE(1)) then
				char1RE <= "-11.8125";
			elsif QstateRE(1) = to_sfixed(-11.7500,QstateRE(1)) then
				char1RE <= "-11.7500";
			elsif QstateRE(1) = to_sfixed(-11.6875,QstateRE(1)) then
				char1RE <= "-11.6875";
			elsif QstateRE(1) = to_sfixed(-11.6250,QstateRE(1)) then
				char1RE <= "-11.6250";
			elsif QstateRE(1) = to_sfixed(-11.5625,QstateRE(1)) then
				char1RE <= "-11.5625";
			elsif QstateRE(1) = to_sfixed(-11.5000,QstateRE(1)) then
				char1RE <= "-11.5000";
			elsif QstateRE(1) = to_sfixed(-11.4375,QstateRE(1)) then
				char1RE <= "-11.4375";
			elsif QstateRE(1) = to_sfixed(-11.3750,QstateRE(1)) then
				char1RE <= "-11.3750";
			elsif QstateRE(1) = to_sfixed(-11.3125,QstateRE(1)) then
				char1RE <= "-11.3125";
			elsif QstateRE(1) = to_sfixed(-11.2500,QstateRE(1)) then
				char1RE <= "-11.2500";
			elsif QstateRE(1) = to_sfixed(-11.1875,QstateRE(1)) then
				char1RE <= "-11.1875";
			elsif QstateRE(1) = to_sfixed(-11.1250,QstateRE(1)) then
				char1RE <= "-11.1250";
			elsif QstateRE(1) = to_sfixed(-11.0625,QstateRE(1)) then
				char1RE <= "-11.0625";
			elsif QstateRE(1) = to_sfixed(-11.0000,QstateRE(1)) then
				char1RE <= "-11.0000";
			elsif QstateRE(1) = to_sfixed(-10.9375,QstateRE(1)) then
				char1RE <= "-10.9375";
			elsif QstateRE(1) = to_sfixed(-10.8750,QstateRE(1)) then
				char1RE <= "-10.8750";
			elsif QstateRE(1) = to_sfixed(-10.8125,QstateRE(1)) then
				char1RE <= "-10.8125";
			elsif QstateRE(1) = to_sfixed(-10.7500,QstateRE(1)) then
				char1RE <= "-10.7500";
			elsif QstateRE(1) = to_sfixed(-10.6875,QstateRE(1)) then
				char1RE <= "-10.6875";
			elsif QstateRE(1) = to_sfixed(-10.6250,QstateRE(1)) then
				char1RE <= "-10.6250";
			elsif QstateRE(1) = to_sfixed(-10.5625,QstateRE(1)) then
				char1RE <= "-10.5625";
			elsif QstateRE(1) = to_sfixed(-10.5000,QstateRE(1)) then
				char1RE <= "-10.5000";
			elsif QstateRE(1) = to_sfixed(-10.4375,QstateRE(1)) then
				char1RE <= "-10.4375";
			elsif QstateRE(1) = to_sfixed(-10.3750,QstateRE(1)) then
				char1RE <= "-10.3750";
			elsif QstateRE(1) = to_sfixed(-10.3125,QstateRE(1)) then
				char1RE <= "-10.3125";
			elsif QstateRE(1) = to_sfixed(-10.2500,QstateRE(1)) then
				char1RE <= "-10.2500";
			elsif QstateRE(1) = to_sfixed(-10.1875,QstateRE(1)) then
				char1RE <= "-10.1875";
			elsif QstateRE(1) = to_sfixed(-10.1250,QstateRE(1)) then
				char1RE <= "-10.1250";
			elsif QstateRE(1) = to_sfixed(-10.0625,QstateRE(1)) then
				char1RE <= "-10.0625";
			elsif QstateRE(1) = to_sfixed(-10.0000,QstateRE(1)) then
				char1RE <= "-10.0000";
			elsif QstateRE(1) = to_sfixed(-9.9375,QstateRE(1)) then
				char1RE <= "--9.9375";
			elsif QstateRE(1) = to_sfixed(-9.8750,QstateRE(1)) then
				char1RE <= "--9.8750";
			elsif QstateRE(1) = to_sfixed(-9.8125,QstateRE(1)) then
				char1RE <= "--9.8125";
			elsif QstateRE(1) = to_sfixed(-9.7500,QstateRE(1)) then
				char1RE <= "--9.7500";
			elsif QstateRE(1) = to_sfixed(-9.6875,QstateRE(1)) then
				char1RE <= "--9.6875";
			elsif QstateRE(1) = to_sfixed(-9.6250,QstateRE(1)) then
				char1RE <= "--9.6250";
			elsif QstateRE(1) = to_sfixed(-9.5625,QstateRE(1)) then
				char1RE <= "--9.5625";
			elsif QstateRE(1) = to_sfixed(-9.5000,QstateRE(1)) then
				char1RE <= "--9.5000";
			elsif QstateRE(1) = to_sfixed(-9.4375,QstateRE(1)) then
				char1RE <= "--9.4375";
			elsif QstateRE(1) = to_sfixed(-9.3750,QstateRE(1)) then
				char1RE <= "--9.3750";
			elsif QstateRE(1) = to_sfixed(-9.3125,QstateRE(1)) then
				char1RE <= "--9.3125";
			elsif QstateRE(1) = to_sfixed(-9.2500,QstateRE(1)) then
				char1RE <= "--9.2500";
			elsif QstateRE(1) = to_sfixed(-9.1875,QstateRE(1)) then
				char1RE <= "--9.1875";
			elsif QstateRE(1) = to_sfixed(-9.1250,QstateRE(1)) then
				char1RE <= "--9.1250";
			elsif QstateRE(1) = to_sfixed(-9.0625,QstateRE(1)) then
				char1RE <= "--9.0625";
			elsif QstateRE(1) = to_sfixed(-9.0000,QstateRE(1)) then
				char1RE <= "--9.0000";
			elsif QstateRE(1) = to_sfixed(-8.9375,QstateRE(1)) then
				char1RE <= "--8.9375";
			elsif QstateRE(1) = to_sfixed(-8.8750,QstateRE(1)) then
				char1RE <= "--8.8750";
			elsif QstateRE(1) = to_sfixed(-8.8125,QstateRE(1)) then
				char1RE <= "--8.8125";
			elsif QstateRE(1) = to_sfixed(-8.7500,QstateRE(1)) then
				char1RE <= "--8.7500";
			elsif QstateRE(1) = to_sfixed(-8.6875,QstateRE(1)) then
				char1RE <= "--8.6875";
			elsif QstateRE(1) = to_sfixed(-8.6250,QstateRE(1)) then
				char1RE <= "--8.6250";
			elsif QstateRE(1) = to_sfixed(-8.5625,QstateRE(1)) then
				char1RE <= "--8.5625";
			elsif QstateRE(1) = to_sfixed(-8.5000,QstateRE(1)) then
				char1RE <= "--8.5000";
			elsif QstateRE(1) = to_sfixed(-8.4375,QstateRE(1)) then
				char1RE <= "--8.4375";
			elsif QstateRE(1) = to_sfixed(-8.3750,QstateRE(1)) then
				char1RE <= "--8.3750";
			elsif QstateRE(1) = to_sfixed(-8.3125,QstateRE(1)) then
				char1RE <= "--8.3125";
			elsif QstateRE(1) = to_sfixed(-8.2500,QstateRE(1)) then
				char1RE <= "--8.2500";
			elsif QstateRE(1) = to_sfixed(-8.1875,QstateRE(1)) then
				char1RE <= "--8.1875";
			elsif QstateRE(1) = to_sfixed(-8.1250,QstateRE(1)) then
				char1RE <= "--8.1250";
			elsif QstateRE(1) = to_sfixed(-8.0625,QstateRE(1)) then
				char1RE <= "--8.0625";
			elsif QstateRE(1) = to_sfixed(-8.0000,QstateRE(1)) then
				char1RE <= "--8.0000";
			elsif QstateRE(1) = to_sfixed(-7.9375,QstateRE(1)) then
				char1RE <= "--7.9375";
			elsif QstateRE(1) = to_sfixed(-7.8750,QstateRE(1)) then
				char1RE <= "--7.8750";
			elsif QstateRE(1) = to_sfixed(-7.8125,QstateRE(1)) then
				char1RE <= "--7.8125";
			elsif QstateRE(1) = to_sfixed(-7.7500,QstateRE(1)) then
				char1RE <= "--7.7500";
			elsif QstateRE(1) = to_sfixed(-7.6875,QstateRE(1)) then
				char1RE <= "--7.6875";
			elsif QstateRE(1) = to_sfixed(-7.6250,QstateRE(1)) then
				char1RE <= "--7.6250";
			elsif QstateRE(1) = to_sfixed(-7.5625,QstateRE(1)) then
				char1RE <= "--7.5625";
			elsif QstateRE(1) = to_sfixed(-7.5000,QstateRE(1)) then
				char1RE <= "--7.5000";
			elsif QstateRE(1) = to_sfixed(-7.4375,QstateRE(1)) then
				char1RE <= "--7.4375";
			elsif QstateRE(1) = to_sfixed(-7.3750,QstateRE(1)) then
				char1RE <= "--7.3750";
			elsif QstateRE(1) = to_sfixed(-7.3125,QstateRE(1)) then
				char1RE <= "--7.3125";
			elsif QstateRE(1) = to_sfixed(-7.2500,QstateRE(1)) then
				char1RE <= "--7.2500";
			elsif QstateRE(1) = to_sfixed(-7.1875,QstateRE(1)) then
				char1RE <= "--7.1875";
			elsif QstateRE(1) = to_sfixed(-7.1250,QstateRE(1)) then
				char1RE <= "--7.1250";
			elsif QstateRE(1) = to_sfixed(-7.0625,QstateRE(1)) then
				char1RE <= "--7.0625";
			elsif QstateRE(1) = to_sfixed(-7.0000,QstateRE(1)) then
				char1RE <= "--7.0000";
			elsif QstateRE(1) = to_sfixed(-6.9375,QstateRE(1)) then
				char1RE <= "--6.9375";
			elsif QstateRE(1) = to_sfixed(-6.8750,QstateRE(1)) then
				char1RE <= "--6.8750";
			elsif QstateRE(1) = to_sfixed(-6.8125,QstateRE(1)) then
				char1RE <= "--6.8125";
			elsif QstateRE(1) = to_sfixed(-6.7500,QstateRE(1)) then
				char1RE <= "--6.7500";
			elsif QstateRE(1) = to_sfixed(-6.6875,QstateRE(1)) then
				char1RE <= "--6.6875";
			elsif QstateRE(1) = to_sfixed(-6.6250,QstateRE(1)) then
				char1RE <= "--6.6250";
			elsif QstateRE(1) = to_sfixed(-6.5625,QstateRE(1)) then
				char1RE <= "--6.5625";
			elsif QstateRE(1) = to_sfixed(-6.5000,QstateRE(1)) then
				char1RE <= "--6.5000";
			elsif QstateRE(1) = to_sfixed(-6.4375,QstateRE(1)) then
				char1RE <= "--6.4375";
			elsif QstateRE(1) = to_sfixed(-6.3750,QstateRE(1)) then
				char1RE <= "--6.3750";
			elsif QstateRE(1) = to_sfixed(-6.3125,QstateRE(1)) then
				char1RE <= "--6.3125";
			elsif QstateRE(1) = to_sfixed(-6.2500,QstateRE(1)) then
				char1RE <= "--6.2500";
			elsif QstateRE(1) = to_sfixed(-6.1875,QstateRE(1)) then
				char1RE <= "--6.1875";
			elsif QstateRE(1) = to_sfixed(-6.1250,QstateRE(1)) then
				char1RE <= "--6.1250";
			elsif QstateRE(1) = to_sfixed(-6.0625,QstateRE(1)) then
				char1RE <= "--6.0625";
			elsif QstateRE(1) = to_sfixed(-6.0000,QstateRE(1)) then
				char1RE <= "--6.0000";
			elsif QstateRE(1) = to_sfixed(-5.9375,QstateRE(1)) then
				char1RE <= "--5.9375";
			elsif QstateRE(1) = to_sfixed(-5.8750,QstateRE(1)) then
				char1RE <= "--5.8750";
			elsif QstateRE(1) = to_sfixed(-5.8125,QstateRE(1)) then
				char1RE <= "--5.8125";
			elsif QstateRE(1) = to_sfixed(-5.7500,QstateRE(1)) then
				char1RE <= "--5.7500";
			elsif QstateRE(1) = to_sfixed(-5.6875,QstateRE(1)) then
				char1RE <= "--5.6875";
			elsif QstateRE(1) = to_sfixed(-5.6250,QstateRE(1)) then
				char1RE <= "--5.6250";
			elsif QstateRE(1) = to_sfixed(-5.5625,QstateRE(1)) then
				char1RE <= "--5.5625";
			elsif QstateRE(1) = to_sfixed(-5.5000,QstateRE(1)) then
				char1RE <= "--5.5000";
			elsif QstateRE(1) = to_sfixed(-5.4375,QstateRE(1)) then
				char1RE <= "--5.4375";
			elsif QstateRE(1) = to_sfixed(-5.3750,QstateRE(1)) then
				char1RE <= "--5.3750";
			elsif QstateRE(1) = to_sfixed(-5.3125,QstateRE(1)) then
				char1RE <= "--5.3125";
			elsif QstateRE(1) = to_sfixed(-5.2500,QstateRE(1)) then
				char1RE <= "--5.2500";
			elsif QstateRE(1) = to_sfixed(-5.1875,QstateRE(1)) then
				char1RE <= "--5.1875";
			elsif QstateRE(1) = to_sfixed(-5.1250,QstateRE(1)) then
				char1RE <= "--5.1250";
			elsif QstateRE(1) = to_sfixed(-5.0625,QstateRE(1)) then
				char1RE <= "--5.0625";
			elsif QstateRE(1) = to_sfixed(-5.0000,QstateRE(1)) then
				char1RE <= "--5.0000";
			elsif QstateRE(1) = to_sfixed(-4.9375,QstateRE(1)) then
				char1RE <= "--4.9375";
			elsif QstateRE(1) = to_sfixed(-4.8750,QstateRE(1)) then
				char1RE <= "--4.8750";
			elsif QstateRE(1) = to_sfixed(-4.8125,QstateRE(1)) then
				char1RE <= "--4.8125";
			elsif QstateRE(1) = to_sfixed(-4.7500,QstateRE(1)) then
				char1RE <= "--4.7500";
			elsif QstateRE(1) = to_sfixed(-4.6875,QstateRE(1)) then
				char1RE <= "--4.6875";
			elsif QstateRE(1) = to_sfixed(-4.6250,QstateRE(1)) then
				char1RE <= "--4.6250";
			elsif QstateRE(1) = to_sfixed(-4.5625,QstateRE(1)) then
				char1RE <= "--4.5625";
			elsif QstateRE(1) = to_sfixed(-4.5000,QstateRE(1)) then
				char1RE <= "--4.5000";
			elsif QstateRE(1) = to_sfixed(-4.4375,QstateRE(1)) then
				char1RE <= "--4.4375";
			elsif QstateRE(1) = to_sfixed(-4.3750,QstateRE(1)) then
				char1RE <= "--4.3750";
			elsif QstateRE(1) = to_sfixed(-4.3125,QstateRE(1)) then
				char1RE <= "--4.3125";
			elsif QstateRE(1) = to_sfixed(-4.2500,QstateRE(1)) then
				char1RE <= "--4.2500";
			elsif QstateRE(1) = to_sfixed(-4.1875,QstateRE(1)) then
				char1RE <= "--4.1875";
			elsif QstateRE(1) = to_sfixed(-4.1250,QstateRE(1)) then
				char1RE <= "--4.1250";
			elsif QstateRE(1) = to_sfixed(-4.0625,QstateRE(1)) then
				char1RE <= "--4.0625";
			elsif QstateRE(1) = to_sfixed(-4.0000,QstateRE(1)) then
				char1RE <= "--4.0000";
			elsif QstateRE(1) = to_sfixed(-3.9375,QstateRE(1)) then
				char1RE <= "--3.9375";
			elsif QstateRE(1) = to_sfixed(-3.8750,QstateRE(1)) then
				char1RE <= "--3.8750";
			elsif QstateRE(1) = to_sfixed(-3.8125,QstateRE(1)) then
				char1RE <= "--3.8125";
			elsif QstateRE(1) = to_sfixed(-3.7500,QstateRE(1)) then
				char1RE <= "--3.7500";
			elsif QstateRE(1) = to_sfixed(-3.6875,QstateRE(1)) then
				char1RE <= "--3.6875";
			elsif QstateRE(1) = to_sfixed(-3.6250,QstateRE(1)) then
				char1RE <= "--3.6250";
			elsif QstateRE(1) = to_sfixed(-3.5625,QstateRE(1)) then
				char1RE <= "--3.5625";
			elsif QstateRE(1) = to_sfixed(-3.5000,QstateRE(1)) then
				char1RE <= "--3.5000";
			elsif QstateRE(1) = to_sfixed(-3.4375,QstateRE(1)) then
				char1RE <= "--3.4375";
			elsif QstateRE(1) = to_sfixed(-3.3750,QstateRE(1)) then
				char1RE <= "--3.3750";
			elsif QstateRE(1) = to_sfixed(-3.3125,QstateRE(1)) then
				char1RE <= "--3.3125";
			elsif QstateRE(1) = to_sfixed(-3.2500,QstateRE(1)) then
				char1RE <= "--3.2500";
			elsif QstateRE(1) = to_sfixed(-3.1875,QstateRE(1)) then
				char1RE <= "--3.1875";
			elsif QstateRE(1) = to_sfixed(-3.1250,QstateRE(1)) then
				char1RE <= "--3.1250";
			elsif QstateRE(1) = to_sfixed(-3.0625,QstateRE(1)) then
				char1RE <= "--3.0625";
			elsif QstateRE(1) = to_sfixed(-3.0000,QstateRE(1)) then
				char1RE <= "--3.0000";
			elsif QstateRE(1) = to_sfixed(-2.9375,QstateRE(1)) then
				char1RE <= "--2.9375";
			elsif QstateRE(1) = to_sfixed(-2.8750,QstateRE(1)) then
				char1RE <= "--2.8750";
			elsif QstateRE(1) = to_sfixed(-2.8125,QstateRE(1)) then
				char1RE <= "--2.8125";
			elsif QstateRE(1) = to_sfixed(-2.7500,QstateRE(1)) then
				char1RE <= "--2.7500";
			elsif QstateRE(1) = to_sfixed(-2.6875,QstateRE(1)) then
				char1RE <= "--2.6875";
			elsif QstateRE(1) = to_sfixed(-2.6250,QstateRE(1)) then
				char1RE <= "--2.6250";
			elsif QstateRE(1) = to_sfixed(-2.5625,QstateRE(1)) then
				char1RE <= "--2.5625";
			elsif QstateRE(1) = to_sfixed(-2.5000,QstateRE(1)) then
				char1RE <= "--2.5000";
			elsif QstateRE(1) = to_sfixed(-2.4375,QstateRE(1)) then
				char1RE <= "--2.4375";
			elsif QstateRE(1) = to_sfixed(-2.3750,QstateRE(1)) then
				char1RE <= "--2.3750";
			elsif QstateRE(1) = to_sfixed(-2.3125,QstateRE(1)) then
				char1RE <= "--2.3125";
			elsif QstateRE(1) = to_sfixed(-2.2500,QstateRE(1)) then
				char1RE <= "--2.2500";
			elsif QstateRE(1) = to_sfixed(-2.1875,QstateRE(1)) then
				char1RE <= "--2.1875";
			elsif QstateRE(1) = to_sfixed(-2.1250,QstateRE(1)) then
				char1RE <= "--2.1250";
			elsif QstateRE(1) = to_sfixed(-2.0625,QstateRE(1)) then
				char1RE <= "--2.0625";
			elsif QstateRE(1) = to_sfixed(-2.0000,QstateRE(1)) then
				char1RE <= "--2.0000";
			elsif QstateRE(1) = to_sfixed(-1.9375,QstateRE(1)) then
				char1RE <= "--1.9375";
			elsif QstateRE(1) = to_sfixed(-1.8750,QstateRE(1)) then
				char1RE <= "--1.8750";
			elsif QstateRE(1) = to_sfixed(-1.8125,QstateRE(1)) then
				char1RE <= "--1.8125";
			elsif QstateRE(1) = to_sfixed(-1.7500,QstateRE(1)) then
				char1RE <= "--1.7500";
			elsif QstateRE(1) = to_sfixed(-1.6875,QstateRE(1)) then
				char1RE <= "--1.6875";
			elsif QstateRE(1) = to_sfixed(-1.6250,QstateRE(1)) then
				char1RE <= "--1.6250";
			elsif QstateRE(1) = to_sfixed(-1.5625,QstateRE(1)) then
				char1RE <= "--1.5625";
			elsif QstateRE(1) = to_sfixed(-1.5000,QstateRE(1)) then
				char1RE <= "--1.5000";
			elsif QstateRE(1) = to_sfixed(-1.4375,QstateRE(1)) then
				char1RE <= "--1.4375";
			elsif QstateRE(1) = to_sfixed(-1.3750,QstateRE(1)) then
				char1RE <= "--1.3750";
			elsif QstateRE(1) = to_sfixed(-1.3125,QstateRE(1)) then
				char1RE <= "--1.3125";
			elsif QstateRE(1) = to_sfixed(-1.2500,QstateRE(1)) then
				char1RE <= "--1.2500";
			elsif QstateRE(1) = to_sfixed(-1.1875,QstateRE(1)) then
				char1RE <= "--1.1875";
			elsif QstateRE(1) = to_sfixed(-1.1250,QstateRE(1)) then
				char1RE <= "--1.1250";
			elsif QstateRE(1) = to_sfixed(-1.0625,QstateRE(1)) then
				char1RE <= "--1.0625";
			elsif QstateRE(1) = to_sfixed(-1.0000,QstateRE(1)) then
				char1RE <= "--1.0000";
			elsif QstateRE(1) = to_sfixed(-0.9375,QstateRE(1)) then
				char1RE <= "--0.9375";
			elsif QstateRE(1) = to_sfixed(-0.8750,QstateRE(1)) then
				char1RE <= "--0.8750";
			elsif QstateRE(1) = to_sfixed(-0.8125,QstateRE(1)) then
				char1RE <= "--0.8125";
			elsif QstateRE(1) = to_sfixed(-0.7500,QstateRE(1)) then
				char1RE <= "--0.7500";
			elsif QstateRE(1) = to_sfixed(-0.6875,QstateRE(1)) then
				char1RE <= "--0.6875";
			elsif QstateRE(1) = to_sfixed(-0.6250,QstateRE(1)) then
				char1RE <= "--0.6250";
			elsif QstateRE(1) = to_sfixed(-0.5625,QstateRE(1)) then
				char1RE <= "--0.5625";
			elsif QstateRE(1) = to_sfixed(-0.5000,QstateRE(1)) then
				char1RE <= "--0.5000";
			elsif QstateRE(1) = to_sfixed(-0.4375,QstateRE(1)) then
				char1RE <= "--0.4375";
			elsif QstateRE(1) = to_sfixed(-0.3750,QstateRE(1)) then
				char1RE <= "--0.3750";
			elsif QstateRE(1) = to_sfixed(-0.3125,QstateRE(1)) then
				char1RE <= "--0.3125";
			elsif QstateRE(1) = to_sfixed(-0.2500,QstateRE(1)) then
				char1RE <= "--0.2500";
			elsif QstateRE(1) = to_sfixed(-0.1875,QstateRE(1)) then
				char1RE <= "--0.1875";
			elsif QstateRE(1) = to_sfixed(-0.1250,QstateRE(1)) then
				char1RE <= "--0.1250";
			elsif QstateRE(1) = to_sfixed(-0.0625,QstateRE(1)) then
				char1RE <= "--0.0625";
			elsif QstateRE(1) = to_sfixed(00.0000,QstateRE(1)) then
				char1RE <= "+00.0000";
			elsif QstateRE(1) = to_sfixed(00.0625,QstateRE(1)) then
				char1RE <= "+00.0625";
			elsif QstateRE(1) = to_sfixed(00.1250,QstateRE(1)) then
				char1RE <= "+00.1250";
			elsif QstateRE(1) = to_sfixed(00.1875,QstateRE(1)) then
				char1RE <= "+00.1875";
			elsif QstateRE(1) = to_sfixed(00.2500,QstateRE(1)) then
				char1RE <= "+00.2500";
			elsif QstateRE(1) = to_sfixed(00.3125,QstateRE(1)) then
				char1RE <= "+00.3125";
			elsif QstateRE(1) = to_sfixed(00.3750,QstateRE(1)) then
				char1RE <= "+00.3750";
			elsif QstateRE(1) = to_sfixed(00.4375,QstateRE(1)) then
				char1RE <= "+00.4375";
			elsif QstateRE(1) = to_sfixed(00.5000,QstateRE(1)) then
				char1RE <= "+00.5000";
			elsif QstateRE(1) = to_sfixed(00.5625,QstateRE(1)) then
				char1RE <= "+00.5625";
			elsif QstateRE(1) = to_sfixed(00.6250,QstateRE(1)) then
				char1RE <= "+00.6250";
			elsif QstateRE(1) = to_sfixed(00.6875,QstateRE(1)) then
				char1RE <= "+00.6875";
			elsif QstateRE(1) = to_sfixed(00.7500,QstateRE(1)) then
				char1RE <= "+00.7500";
			elsif QstateRE(1) = to_sfixed(00.8125,QstateRE(1)) then
				char1RE <= "+00.8125";
			elsif QstateRE(1) = to_sfixed(00.8750,QstateRE(1)) then
				char1RE <= "+00.8750";
			elsif QstateRE(1) = to_sfixed(00.9375,QstateRE(1)) then
				char1RE <= "+00.9375";
			elsif QstateRE(1) = to_sfixed(01.0000,QstateRE(1)) then
				char1RE <= "+01.0000";
			elsif QstateRE(1) = to_sfixed(01.0625,QstateRE(1)) then
				char1RE <= "+01.0625";
			elsif QstateRE(1) = to_sfixed(01.1250,QstateRE(1)) then
				char1RE <= "+01.1250";
			elsif QstateRE(1) = to_sfixed(01.1875,QstateRE(1)) then
				char1RE <= "+01.1875";
			elsif QstateRE(1) = to_sfixed(01.2500,QstateRE(1)) then
				char1RE <= "+01.2500";
			elsif QstateRE(1) = to_sfixed(01.3125,QstateRE(1)) then
				char1RE <= "+01.3125";
			elsif QstateRE(1) = to_sfixed(01.3750,QstateRE(1)) then
				char1RE <= "+01.3750";
			elsif QstateRE(1) = to_sfixed(01.4375,QstateRE(1)) then
				char1RE <= "+01.4375";
			elsif QstateRE(1) = to_sfixed(01.5000,QstateRE(1)) then
				char1RE <= "+01.5000";
			elsif QstateRE(1) = to_sfixed(01.5625,QstateRE(1)) then
				char1RE <= "+01.5625";
			elsif QstateRE(1) = to_sfixed(01.6250,QstateRE(1)) then
				char1RE <= "+01.6250";
			elsif QstateRE(1) = to_sfixed(01.6875,QstateRE(1)) then
				char1RE <= "+01.6875";
			elsif QstateRE(1) = to_sfixed(01.7500,QstateRE(1)) then
				char1RE <= "+01.7500";
			elsif QstateRE(1) = to_sfixed(01.8125,QstateRE(1)) then
				char1RE <= "+01.8125";
			elsif QstateRE(1) = to_sfixed(01.8750,QstateRE(1)) then
				char1RE <= "+01.8750";
			elsif QstateRE(1) = to_sfixed(01.9375,QstateRE(1)) then
				char1RE <= "+01.9375";
			elsif QstateRE(1) = to_sfixed(02.0000,QstateRE(1)) then
				char1RE <= "+02.0000";
			elsif QstateRE(1) = to_sfixed(02.0625,QstateRE(1)) then
				char1RE <= "+02.0625";
			elsif QstateRE(1) = to_sfixed(02.1250,QstateRE(1)) then
				char1RE <= "+02.1250";
			elsif QstateRE(1) = to_sfixed(02.1875,QstateRE(1)) then
				char1RE <= "+02.1875";
			elsif QstateRE(1) = to_sfixed(02.2500,QstateRE(1)) then
				char1RE <= "+02.2500";
			elsif QstateRE(1) = to_sfixed(02.3125,QstateRE(1)) then
				char1RE <= "+02.3125";
			elsif QstateRE(1) = to_sfixed(02.3750,QstateRE(1)) then
				char1RE <= "+02.3750";
			elsif QstateRE(1) = to_sfixed(02.4375,QstateRE(1)) then
				char1RE <= "+02.4375";
			elsif QstateRE(1) = to_sfixed(02.5000,QstateRE(1)) then
				char1RE <= "+02.5000";
			elsif QstateRE(1) = to_sfixed(02.5625,QstateRE(1)) then
				char1RE <= "+02.5625";
			elsif QstateRE(1) = to_sfixed(02.6250,QstateRE(1)) then
				char1RE <= "+02.6250";
			elsif QstateRE(1) = to_sfixed(02.6875,QstateRE(1)) then
				char1RE <= "+02.6875";
			elsif QstateRE(1) = to_sfixed(02.7500,QstateRE(1)) then
				char1RE <= "+02.7500";
			elsif QstateRE(1) = to_sfixed(02.8125,QstateRE(1)) then
				char1RE <= "+02.8125";
			elsif QstateRE(1) = to_sfixed(02.8750,QstateRE(1)) then
				char1RE <= "+02.8750";
			elsif QstateRE(1) = to_sfixed(02.9375,QstateRE(1)) then
				char1RE <= "+02.9375";
			elsif QstateRE(1) = to_sfixed(03.0000,QstateRE(1)) then
				char1RE <= "+03.0000";
			elsif QstateRE(1) = to_sfixed(03.0625,QstateRE(1)) then
				char1RE <= "+03.0625";
			elsif QstateRE(1) = to_sfixed(03.1250,QstateRE(1)) then
				char1RE <= "+03.1250";
			elsif QstateRE(1) = to_sfixed(03.1875,QstateRE(1)) then
				char1RE <= "+03.1875";
			elsif QstateRE(1) = to_sfixed(03.2500,QstateRE(1)) then
				char1RE <= "+03.2500";
			elsif QstateRE(1) = to_sfixed(03.3125,QstateRE(1)) then
				char1RE <= "+03.3125";
			elsif QstateRE(1) = to_sfixed(03.3750,QstateRE(1)) then
				char1RE <= "+03.3750";
			elsif QstateRE(1) = to_sfixed(03.4375,QstateRE(1)) then
				char1RE <= "+03.4375";
			elsif QstateRE(1) = to_sfixed(03.5000,QstateRE(1)) then
				char1RE <= "+03.5000";
			elsif QstateRE(1) = to_sfixed(03.5625,QstateRE(1)) then
				char1RE <= "+03.5625";
			elsif QstateRE(1) = to_sfixed(03.6250,QstateRE(1)) then
				char1RE <= "+03.6250";
			elsif QstateRE(1) = to_sfixed(03.6875,QstateRE(1)) then
				char1RE <= "+03.6875";
			elsif QstateRE(1) = to_sfixed(03.7500,QstateRE(1)) then
				char1RE <= "+03.7500";
			elsif QstateRE(1) = to_sfixed(03.8125,QstateRE(1)) then
				char1RE <= "+03.8125";
			elsif QstateRE(1) = to_sfixed(03.8750,QstateRE(1)) then
				char1RE <= "+03.8750";
			elsif QstateRE(1) = to_sfixed(03.9375,QstateRE(1)) then
				char1RE <= "+03.9375";
			elsif QstateRE(1) = to_sfixed(04.0000,QstateRE(1)) then
				char1RE <= "+04.0000";
			elsif QstateRE(1) = to_sfixed(04.0625,QstateRE(1)) then
				char1RE <= "+04.0625";
			elsif QstateRE(1) = to_sfixed(04.1250,QstateRE(1)) then
				char1RE <= "+04.1250";
			elsif QstateRE(1) = to_sfixed(04.1875,QstateRE(1)) then
				char1RE <= "+04.1875";
			elsif QstateRE(1) = to_sfixed(04.2500,QstateRE(1)) then
				char1RE <= "+04.2500";
			elsif QstateRE(1) = to_sfixed(04.3125,QstateRE(1)) then
				char1RE <= "+04.3125";
			elsif QstateRE(1) = to_sfixed(04.3750,QstateRE(1)) then
				char1RE <= "+04.3750";
			elsif QstateRE(1) = to_sfixed(04.4375,QstateRE(1)) then
				char1RE <= "+04.4375";
			elsif QstateRE(1) = to_sfixed(04.5000,QstateRE(1)) then
				char1RE <= "+04.5000";
			elsif QstateRE(1) = to_sfixed(04.5625,QstateRE(1)) then
				char1RE <= "+04.5625";
			elsif QstateRE(1) = to_sfixed(04.6250,QstateRE(1)) then
				char1RE <= "+04.6250";
			elsif QstateRE(1) = to_sfixed(04.6875,QstateRE(1)) then
				char1RE <= "+04.6875";
			elsif QstateRE(1) = to_sfixed(04.7500,QstateRE(1)) then
				char1RE <= "+04.7500";
			elsif QstateRE(1) = to_sfixed(04.8125,QstateRE(1)) then
				char1RE <= "+04.8125";
			elsif QstateRE(1) = to_sfixed(04.8750,QstateRE(1)) then
				char1RE <= "+04.8750";
			elsif QstateRE(1) = to_sfixed(04.9375,QstateRE(1)) then
				char1RE <= "+04.9375";
			elsif QstateRE(1) = to_sfixed(05.0000,QstateRE(1)) then
				char1RE <= "+05.0000";
			elsif QstateRE(1) = to_sfixed(05.0625,QstateRE(1)) then
				char1RE <= "+05.0625";
			elsif QstateRE(1) = to_sfixed(05.1250,QstateRE(1)) then
				char1RE <= "+05.1250";
			elsif QstateRE(1) = to_sfixed(05.1875,QstateRE(1)) then
				char1RE <= "+05.1875";
			elsif QstateRE(1) = to_sfixed(05.2500,QstateRE(1)) then
				char1RE <= "+05.2500";
			elsif QstateRE(1) = to_sfixed(05.3125,QstateRE(1)) then
				char1RE <= "+05.3125";
			elsif QstateRE(1) = to_sfixed(05.3750,QstateRE(1)) then
				char1RE <= "+05.3750";
			elsif QstateRE(1) = to_sfixed(05.4375,QstateRE(1)) then
				char1RE <= "+05.4375";
			elsif QstateRE(1) = to_sfixed(05.5000,QstateRE(1)) then
				char1RE <= "+05.5000";
			elsif QstateRE(1) = to_sfixed(05.5625,QstateRE(1)) then
				char1RE <= "+05.5625";
			elsif QstateRE(1) = to_sfixed(05.6250,QstateRE(1)) then
				char1RE <= "+05.6250";
			elsif QstateRE(1) = to_sfixed(05.6875,QstateRE(1)) then
				char1RE <= "+05.6875";
			elsif QstateRE(1) = to_sfixed(05.7500,QstateRE(1)) then
				char1RE <= "+05.7500";
			elsif QstateRE(1) = to_sfixed(05.8125,QstateRE(1)) then
				char1RE <= "+05.8125";
			elsif QstateRE(1) = to_sfixed(05.8750,QstateRE(1)) then
				char1RE <= "+05.8750";
			elsif QstateRE(1) = to_sfixed(05.9375,QstateRE(1)) then
				char1RE <= "+05.9375";
			elsif QstateRE(1) = to_sfixed(06.0000,QstateRE(1)) then
				char1RE <= "+06.0000";
			elsif QstateRE(1) = to_sfixed(06.0625,QstateRE(1)) then
				char1RE <= "+06.0625";
			elsif QstateRE(1) = to_sfixed(06.1250,QstateRE(1)) then
				char1RE <= "+06.1250";
			elsif QstateRE(1) = to_sfixed(06.1875,QstateRE(1)) then
				char1RE <= "+06.1875";
			elsif QstateRE(1) = to_sfixed(06.2500,QstateRE(1)) then
				char1RE <= "+06.2500";
			elsif QstateRE(1) = to_sfixed(06.3125,QstateRE(1)) then
				char1RE <= "+06.3125";
			elsif QstateRE(1) = to_sfixed(06.3750,QstateRE(1)) then
				char1RE <= "+06.3750";
			elsif QstateRE(1) = to_sfixed(06.4375,QstateRE(1)) then
				char1RE <= "+06.4375";
			elsif QstateRE(1) = to_sfixed(06.5000,QstateRE(1)) then
				char1RE <= "+06.5000";
			elsif QstateRE(1) = to_sfixed(06.5625,QstateRE(1)) then
				char1RE <= "+06.5625";
			elsif QstateRE(1) = to_sfixed(06.6250,QstateRE(1)) then
				char1RE <= "+06.6250";
			elsif QstateRE(1) = to_sfixed(06.6875,QstateRE(1)) then
				char1RE <= "+06.6875";
			elsif QstateRE(1) = to_sfixed(06.7500,QstateRE(1)) then
				char1RE <= "+06.7500";
			elsif QstateRE(1) = to_sfixed(06.8125,QstateRE(1)) then
				char1RE <= "+06.8125";
			elsif QstateRE(1) = to_sfixed(06.8750,QstateRE(1)) then
				char1RE <= "+06.8750";
			elsif QstateRE(1) = to_sfixed(06.9375,QstateRE(1)) then
				char1RE <= "+06.9375";
			elsif QstateRE(1) = to_sfixed(07.0000,QstateRE(1)) then
				char1RE <= "+07.0000";
			elsif QstateRE(1) = to_sfixed(07.0625,QstateRE(1)) then
				char1RE <= "+07.0625";
			elsif QstateRE(1) = to_sfixed(07.1250,QstateRE(1)) then
				char1RE <= "+07.1250";
			elsif QstateRE(1) = to_sfixed(07.1875,QstateRE(1)) then
				char1RE <= "+07.1875";
			elsif QstateRE(1) = to_sfixed(07.2500,QstateRE(1)) then
				char1RE <= "+07.2500";
			elsif QstateRE(1) = to_sfixed(07.3125,QstateRE(1)) then
				char1RE <= "+07.3125";
			elsif QstateRE(1) = to_sfixed(07.3750,QstateRE(1)) then
				char1RE <= "+07.3750";
			elsif QstateRE(1) = to_sfixed(07.4375,QstateRE(1)) then
				char1RE <= "+07.4375";
			elsif QstateRE(1) = to_sfixed(07.5000,QstateRE(1)) then
				char1RE <= "+07.5000";
			elsif QstateRE(1) = to_sfixed(07.5625,QstateRE(1)) then
				char1RE <= "+07.5625";
			elsif QstateRE(1) = to_sfixed(07.6250,QstateRE(1)) then
				char1RE <= "+07.6250";
			elsif QstateRE(1) = to_sfixed(07.6875,QstateRE(1)) then
				char1RE <= "+07.6875";
			elsif QstateRE(1) = to_sfixed(07.7500,QstateRE(1)) then
				char1RE <= "+07.7500";
			elsif QstateRE(1) = to_sfixed(07.8125,QstateRE(1)) then
				char1RE <= "+07.8125";
			elsif QstateRE(1) = to_sfixed(07.8750,QstateRE(1)) then
				char1RE <= "+07.8750";
			elsif QstateRE(1) = to_sfixed(07.9375,QstateRE(1)) then
				char1RE <= "+07.9375";
			elsif QstateRE(1) = to_sfixed(08.0000,QstateRE(1)) then
				char1RE <= "+08.0000";
			elsif QstateRE(1) = to_sfixed(08.0625,QstateRE(1)) then
				char1RE <= "+08.0625";
			elsif QstateRE(1) = to_sfixed(08.1250,QstateRE(1)) then
				char1RE <= "+08.1250";
			elsif QstateRE(1) = to_sfixed(08.1875,QstateRE(1)) then
				char1RE <= "+08.1875";
			elsif QstateRE(1) = to_sfixed(08.2500,QstateRE(1)) then
				char1RE <= "+08.2500";
			elsif QstateRE(1) = to_sfixed(08.3125,QstateRE(1)) then
				char1RE <= "+08.3125";
			elsif QstateRE(1) = to_sfixed(08.3750,QstateRE(1)) then
				char1RE <= "+08.3750";
			elsif QstateRE(1) = to_sfixed(08.4375,QstateRE(1)) then
				char1RE <= "+08.4375";
			elsif QstateRE(1) = to_sfixed(08.5000,QstateRE(1)) then
				char1RE <= "+08.5000";
			elsif QstateRE(1) = to_sfixed(08.5625,QstateRE(1)) then
				char1RE <= "+08.5625";
			elsif QstateRE(1) = to_sfixed(08.6250,QstateRE(1)) then
				char1RE <= "+08.6250";
			elsif QstateRE(1) = to_sfixed(08.6875,QstateRE(1)) then
				char1RE <= "+08.6875";
			elsif QstateRE(1) = to_sfixed(08.7500,QstateRE(1)) then
				char1RE <= "+08.7500";
			elsif QstateRE(1) = to_sfixed(08.8125,QstateRE(1)) then
				char1RE <= "+08.8125";
			elsif QstateRE(1) = to_sfixed(08.8750,QstateRE(1)) then
				char1RE <= "+08.8750";
			elsif QstateRE(1) = to_sfixed(08.9375,QstateRE(1)) then
				char1RE <= "+08.9375";
			elsif QstateRE(1) = to_sfixed(09.0000,QstateRE(1)) then
				char1RE <= "+09.0000";
			elsif QstateRE(1) = to_sfixed(09.0625,QstateRE(1)) then
				char1RE <= "+09.0625";
			elsif QstateRE(1) = to_sfixed(09.1250,QstateRE(1)) then
				char1RE <= "+09.1250";
			elsif QstateRE(1) = to_sfixed(09.1875,QstateRE(1)) then
				char1RE <= "+09.1875";
			elsif QstateRE(1) = to_sfixed(09.2500,QstateRE(1)) then
				char1RE <= "+09.2500";
			elsif QstateRE(1) = to_sfixed(09.3125,QstateRE(1)) then
				char1RE <= "+09.3125";
			elsif QstateRE(1) = to_sfixed(09.3750,QstateRE(1)) then
				char1RE <= "+09.3750";
			elsif QstateRE(1) = to_sfixed(09.4375,QstateRE(1)) then
				char1RE <= "+09.4375";
			elsif QstateRE(1) = to_sfixed(09.5000,QstateRE(1)) then
				char1RE <= "+09.5000";
			elsif QstateRE(1) = to_sfixed(09.5625,QstateRE(1)) then
				char1RE <= "+09.5625";
			elsif QstateRE(1) = to_sfixed(09.6250,QstateRE(1)) then
				char1RE <= "+09.6250";
			elsif QstateRE(1) = to_sfixed(09.6875,QstateRE(1)) then
				char1RE <= "+09.6875";
			elsif QstateRE(1) = to_sfixed(09.7500,QstateRE(1)) then
				char1RE <= "+09.7500";
			elsif QstateRE(1) = to_sfixed(09.8125,QstateRE(1)) then
				char1RE <= "+09.8125";
			elsif QstateRE(1) = to_sfixed(09.8750,QstateRE(1)) then
				char1RE <= "+09.8750";
			elsif QstateRE(1) = to_sfixed(09.9375,QstateRE(1)) then
				char1RE <= "+09.9375";
			elsif QstateRE(1) = to_sfixed(10.0000,QstateRE(1)) then
				char1RE <= "+10.0000";
			elsif QstateRE(1) = to_sfixed(10.0625,QstateRE(1)) then
				char1RE <= "+10.0625";
			elsif QstateRE(1) = to_sfixed(10.1250,QstateRE(1)) then
				char1RE <= "+10.1250";
			elsif QstateRE(1) = to_sfixed(10.1875,QstateRE(1)) then
				char1RE <= "+10.1875";
			elsif QstateRE(1) = to_sfixed(10.2500,QstateRE(1)) then
				char1RE <= "+10.2500";
			elsif QstateRE(1) = to_sfixed(10.3125,QstateRE(1)) then
				char1RE <= "+10.3125";
			elsif QstateRE(1) = to_sfixed(10.3750,QstateRE(1)) then
				char1RE <= "+10.3750";
			elsif QstateRE(1) = to_sfixed(10.4375,QstateRE(1)) then
				char1RE <= "+10.4375";
			elsif QstateRE(1) = to_sfixed(10.5000,QstateRE(1)) then
				char1RE <= "+10.5000";
			elsif QstateRE(1) = to_sfixed(10.5625,QstateRE(1)) then
				char1RE <= "+10.5625";
			elsif QstateRE(1) = to_sfixed(10.6250,QstateRE(1)) then
				char1RE <= "+10.6250";
			elsif QstateRE(1) = to_sfixed(10.6875,QstateRE(1)) then
				char1RE <= "+10.6875";
			elsif QstateRE(1) = to_sfixed(10.7500,QstateRE(1)) then
				char1RE <= "+10.7500";
			elsif QstateRE(1) = to_sfixed(10.8125,QstateRE(1)) then
				char1RE <= "+10.8125";
			elsif QstateRE(1) = to_sfixed(10.8750,QstateRE(1)) then
				char1RE <= "+10.8750";
			elsif QstateRE(1) = to_sfixed(10.9375,QstateRE(1)) then
				char1RE <= "+10.9375";
			elsif QstateRE(1) = to_sfixed(11.0000,QstateRE(1)) then
				char1RE <= "+11.0000";
			elsif QstateRE(1) = to_sfixed(11.0625,QstateRE(1)) then
				char1RE <= "+11.0625";
			elsif QstateRE(1) = to_sfixed(11.1250,QstateRE(1)) then
				char1RE <= "+11.1250";
			elsif QstateRE(1) = to_sfixed(11.1875,QstateRE(1)) then
				char1RE <= "+11.1875";
			elsif QstateRE(1) = to_sfixed(11.2500,QstateRE(1)) then
				char1RE <= "+11.2500";
			elsif QstateRE(1) = to_sfixed(11.3125,QstateRE(1)) then
				char1RE <= "+11.3125";
			elsif QstateRE(1) = to_sfixed(11.3750,QstateRE(1)) then
				char1RE <= "+11.3750";
			elsif QstateRE(1) = to_sfixed(11.4375,QstateRE(1)) then
				char1RE <= "+11.4375";
			elsif QstateRE(1) = to_sfixed(11.5000,QstateRE(1)) then
				char1RE <= "+11.5000";
			elsif QstateRE(1) = to_sfixed(11.5625,QstateRE(1)) then
				char1RE <= "+11.5625";
			elsif QstateRE(1) = to_sfixed(11.6250,QstateRE(1)) then
				char1RE <= "+11.6250";
			elsif QstateRE(1) = to_sfixed(11.6875,QstateRE(1)) then
				char1RE <= "+11.6875";
			elsif QstateRE(1) = to_sfixed(11.7500,QstateRE(1)) then
				char1RE <= "+11.7500";
			elsif QstateRE(1) = to_sfixed(11.8125,QstateRE(1)) then
				char1RE <= "+11.8125";
			elsif QstateRE(1) = to_sfixed(11.8750,QstateRE(1)) then
				char1RE <= "+11.8750";
			elsif QstateRE(1) = to_sfixed(11.9375,QstateRE(1)) then
				char1RE <= "+11.9375";
			elsif QstateRE(1) = to_sfixed(12.0000,QstateRE(1)) then
				char1RE <= "+12.0000";
			elsif QstateRE(1) = to_sfixed(12.0625,QstateRE(1)) then
				char1RE <= "+12.0625";
			elsif QstateRE(1) = to_sfixed(12.1250,QstateRE(1)) then
				char1RE <= "+12.1250";
			elsif QstateRE(1) = to_sfixed(12.1875,QstateRE(1)) then
				char1RE <= "+12.1875";
			elsif QstateRE(1) = to_sfixed(12.2500,QstateRE(1)) then
				char1RE <= "+12.2500";
			elsif QstateRE(1) = to_sfixed(12.3125,QstateRE(1)) then
				char1RE <= "+12.3125";
			elsif QstateRE(1) = to_sfixed(12.3750,QstateRE(1)) then
				char1RE <= "+12.3750";
			elsif QstateRE(1) = to_sfixed(12.4375,QstateRE(1)) then
				char1RE <= "+12.4375";
			elsif QstateRE(1) = to_sfixed(12.5000,QstateRE(1)) then
				char1RE <= "+12.5000";
			elsif QstateRE(1) = to_sfixed(12.5625,QstateRE(1)) then
				char1RE <= "+12.5625";
			elsif QstateRE(1) = to_sfixed(12.6250,QstateRE(1)) then
				char1RE <= "+12.6250";
			elsif QstateRE(1) = to_sfixed(12.6875,QstateRE(1)) then
				char1RE <= "+12.6875";
			elsif QstateRE(1) = to_sfixed(12.7500,QstateRE(1)) then
				char1RE <= "+12.7500";
			elsif QstateRE(1) = to_sfixed(12.8125,QstateRE(1)) then
				char1RE <= "+12.8125";
			elsif QstateRE(1) = to_sfixed(12.8750,QstateRE(1)) then
				char1RE <= "+12.8750";
			elsif QstateRE(1) = to_sfixed(12.9375,QstateRE(1)) then
				char1RE <= "+12.9375";
			elsif QstateRE(1) = to_sfixed(13.0000,QstateRE(1)) then
				char1RE <= "+13.0000";
			elsif QstateRE(1) = to_sfixed(13.0625,QstateRE(1)) then
				char1RE <= "+13.0625";
			elsif QstateRE(1) = to_sfixed(13.1250,QstateRE(1)) then
				char1RE <= "+13.1250";
			elsif QstateRE(1) = to_sfixed(13.1875,QstateRE(1)) then
				char1RE <= "+13.1875";
			elsif QstateRE(1) = to_sfixed(13.2500,QstateRE(1)) then
				char1RE <= "+13.2500";
			elsif QstateRE(1) = to_sfixed(13.3125,QstateRE(1)) then
				char1RE <= "+13.3125";
			elsif QstateRE(1) = to_sfixed(13.3750,QstateRE(1)) then
				char1RE <= "+13.3750";
			elsif QstateRE(1) = to_sfixed(13.4375,QstateRE(1)) then
				char1RE <= "+13.4375";
			elsif QstateRE(1) = to_sfixed(13.5000,QstateRE(1)) then
				char1RE <= "+13.5000";
			elsif QstateRE(1) = to_sfixed(13.5625,QstateRE(1)) then
				char1RE <= "+13.5625";
			elsif QstateRE(1) = to_sfixed(13.6250,QstateRE(1)) then
				char1RE <= "+13.6250";
			elsif QstateRE(1) = to_sfixed(13.6875,QstateRE(1)) then
				char1RE <= "+13.6875";
			elsif QstateRE(1) = to_sfixed(13.7500,QstateRE(1)) then
				char1RE <= "+13.7500";
			elsif QstateRE(1) = to_sfixed(13.8125,QstateRE(1)) then
				char1RE <= "+13.8125";
			elsif QstateRE(1) = to_sfixed(13.8750,QstateRE(1)) then
				char1RE <= "+13.8750";
			elsif QstateRE(1) = to_sfixed(13.9375,QstateRE(1)) then
				char1RE <= "+13.9375";
			elsif QstateRE(1) = to_sfixed(14.0000,QstateRE(1)) then
				char1RE <= "+14.0000";
			elsif QstateRE(1) = to_sfixed(14.0625,QstateRE(1)) then
				char1RE <= "+14.0625";
			elsif QstateRE(1) = to_sfixed(14.1250,QstateRE(1)) then
				char1RE <= "+14.1250";
			elsif QstateRE(1) = to_sfixed(14.1875,QstateRE(1)) then
				char1RE <= "+14.1875";
			elsif QstateRE(1) = to_sfixed(14.2500,QstateRE(1)) then
				char1RE <= "+14.2500";
			elsif QstateRE(1) = to_sfixed(14.3125,QstateRE(1)) then
				char1RE <= "+14.3125";
			elsif QstateRE(1) = to_sfixed(14.3750,QstateRE(1)) then
				char1RE <= "+14.3750";
			elsif QstateRE(1) = to_sfixed(14.4375,QstateRE(1)) then
				char1RE <= "+14.4375";
			elsif QstateRE(1) = to_sfixed(14.5000,QstateRE(1)) then
				char1RE <= "+14.5000";
			elsif QstateRE(1) = to_sfixed(14.5625,QstateRE(1)) then
				char1RE <= "+14.5625";
			elsif QstateRE(1) = to_sfixed(14.6250,QstateRE(1)) then
				char1RE <= "+14.6250";
			elsif QstateRE(1) = to_sfixed(14.6875,QstateRE(1)) then
				char1RE <= "+14.6875";
			elsif QstateRE(1) = to_sfixed(14.7500,QstateRE(1)) then
				char1RE <= "+14.7500";
			elsif QstateRE(1) = to_sfixed(14.8125,QstateRE(1)) then
				char1RE <= "+14.8125";
			elsif QstateRE(1) = to_sfixed(14.8750,QstateRE(1)) then
				char1RE <= "+14.8750";
			elsif QstateRE(1) = to_sfixed(14.9375,QstateRE(1)) then
				char1RE <= "+14.9375";
			elsif QstateRE(1) = to_sfixed(15.0000,QstateRE(1)) then
				char1RE <= "+15.0000";
			elsif QstateRE(1) = to_sfixed(15.0625,QstateRE(1)) then
				char1RE <= "+15.0625";
			elsif QstateRE(1) = to_sfixed(15.1250,QstateRE(1)) then
				char1RE <= "+15.1250";
			elsif QstateRE(1) = to_sfixed(15.1875,QstateRE(1)) then
				char1RE <= "+15.1875";
			elsif QstateRE(1) = to_sfixed(15.2500,QstateRE(1)) then
				char1RE <= "+15.2500";
			elsif QstateRE(1) = to_sfixed(15.3125,QstateRE(1)) then
				char1RE <= "+15.3125";
			elsif QstateRE(1) = to_sfixed(15.3750,QstateRE(1)) then
				char1RE <= "+15.3750";
			elsif QstateRE(1) = to_sfixed(15.4375,QstateRE(1)) then
				char1RE <= "+15.4375";
			elsif QstateRE(1) = to_sfixed(15.5000,QstateRE(1)) then
				char1RE <= "+15.5000";
			elsif QstateRE(1) = to_sfixed(15.5625,QstateRE(1)) then
				char1RE <= "+15.5625";
			elsif QstateRE(1) = to_sfixed(15.6250,QstateRE(1)) then
				char1RE <= "+15.6250";
			elsif QstateRE(1) = to_sfixed(15.6875,QstateRE(1)) then
				char1RE <= "+15.6875";
			elsif QstateRE(1) = to_sfixed(15.7500,QstateRE(1)) then
				char1RE <= "+15.7500";
			elsif QstateRE(1) = to_sfixed(15.8125,QstateRE(1)) then
				char1RE <= "+15.8125";
			elsif QstateRE(1) = to_sfixed(15.8750,QstateRE(1)) then
				char1RE <= "+15.8750";
			elsif QstateRE(1) = to_sfixed(15.9375,QstateRE(1)) then
				char1RE <= "+15.9375";
			end if;
			if QstateIM(1) = to_sfixed(-15.9375,QstateIM(1)) then
				char1IM <= "-15.9375";
			elsif QstateIM(1) = to_sfixed(-15.8750,QstateIM(1)) then
				char1IM <= "-15.8750";
			elsif QstateIM(1) = to_sfixed(-15.8125,QstateIM(1)) then
				char1IM <= "-15.8125";
			elsif QstateIM(1) = to_sfixed(-15.7500,QstateIM(1)) then
				char1IM <= "-15.7500";
			elsif QstateIM(1) = to_sfixed(-15.6875,QstateIM(1)) then
				char1IM <= "-15.6875";
			elsif QstateIM(1) = to_sfixed(-15.6250,QstateIM(1)) then
				char1IM <= "-15.6250";
			elsif QstateIM(1) = to_sfixed(-15.5625,QstateIM(1)) then
				char1IM <= "-15.5625";
			elsif QstateIM(1) = to_sfixed(-15.5000,QstateIM(1)) then
				char1IM <= "-15.5000";
			elsif QstateIM(1) = to_sfixed(-15.4375,QstateIM(1)) then
				char1IM <= "-15.4375";
			elsif QstateIM(1) = to_sfixed(-15.3750,QstateIM(1)) then
				char1IM <= "-15.3750";
			elsif QstateIM(1) = to_sfixed(-15.3125,QstateIM(1)) then
				char1IM <= "-15.3125";
			elsif QstateIM(1) = to_sfixed(-15.2500,QstateIM(1)) then
				char1IM <= "-15.2500";
			elsif QstateIM(1) = to_sfixed(-15.1875,QstateIM(1)) then
				char1IM <= "-15.1875";
			elsif QstateIM(1) = to_sfixed(-15.1250,QstateIM(1)) then
				char1IM <= "-15.1250";
			elsif QstateIM(1) = to_sfixed(-15.0625,QstateIM(1)) then
				char1IM <= "-15.0625";
			elsif QstateIM(1) = to_sfixed(-15.0000,QstateIM(1)) then
				char1IM <= "-15.0000";
			elsif QstateIM(1) = to_sfixed(-14.9375,QstateIM(1)) then
				char1IM <= "-14.9375";
			elsif QstateIM(1) = to_sfixed(-14.8750,QstateIM(1)) then
				char1IM <= "-14.8750";
			elsif QstateIM(1) = to_sfixed(-14.8125,QstateIM(1)) then
				char1IM <= "-14.8125";
			elsif QstateIM(1) = to_sfixed(-14.7500,QstateIM(1)) then
				char1IM <= "-14.7500";
			elsif QstateIM(1) = to_sfixed(-14.6875,QstateIM(1)) then
				char1IM <= "-14.6875";
			elsif QstateIM(1) = to_sfixed(-14.6250,QstateIM(1)) then
				char1IM <= "-14.6250";
			elsif QstateIM(1) = to_sfixed(-14.5625,QstateIM(1)) then
				char1IM <= "-14.5625";
			elsif QstateIM(1) = to_sfixed(-14.5000,QstateIM(1)) then
				char1IM <= "-14.5000";
			elsif QstateIM(1) = to_sfixed(-14.4375,QstateIM(1)) then
				char1IM <= "-14.4375";
			elsif QstateIM(1) = to_sfixed(-14.3750,QstateIM(1)) then
				char1IM <= "-14.3750";
			elsif QstateIM(1) = to_sfixed(-14.3125,QstateIM(1)) then
				char1IM <= "-14.3125";
			elsif QstateIM(1) = to_sfixed(-14.2500,QstateIM(1)) then
				char1IM <= "-14.2500";
			elsif QstateIM(1) = to_sfixed(-14.1875,QstateIM(1)) then
				char1IM <= "-14.1875";
			elsif QstateIM(1) = to_sfixed(-14.1250,QstateIM(1)) then
				char1IM <= "-14.1250";
			elsif QstateIM(1) = to_sfixed(-14.0625,QstateIM(1)) then
				char1IM <= "-14.0625";
			elsif QstateIM(1) = to_sfixed(-14.0000,QstateIM(1)) then
				char1IM <= "-14.0000";
			elsif QstateIM(1) = to_sfixed(-13.9375,QstateIM(1)) then
				char1IM <= "-13.9375";
			elsif QstateIM(1) = to_sfixed(-13.8750,QstateIM(1)) then
				char1IM <= "-13.8750";
			elsif QstateIM(1) = to_sfixed(-13.8125,QstateIM(1)) then
				char1IM <= "-13.8125";
			elsif QstateIM(1) = to_sfixed(-13.7500,QstateIM(1)) then
				char1IM <= "-13.7500";
			elsif QstateIM(1) = to_sfixed(-13.6875,QstateIM(1)) then
				char1IM <= "-13.6875";
			elsif QstateIM(1) = to_sfixed(-13.6250,QstateIM(1)) then
				char1IM <= "-13.6250";
			elsif QstateIM(1) = to_sfixed(-13.5625,QstateIM(1)) then
				char1IM <= "-13.5625";
			elsif QstateIM(1) = to_sfixed(-13.5000,QstateIM(1)) then
				char1IM <= "-13.5000";
			elsif QstateIM(1) = to_sfixed(-13.4375,QstateIM(1)) then
				char1IM <= "-13.4375";
			elsif QstateIM(1) = to_sfixed(-13.3750,QstateIM(1)) then
				char1IM <= "-13.3750";
			elsif QstateIM(1) = to_sfixed(-13.3125,QstateIM(1)) then
				char1IM <= "-13.3125";
			elsif QstateIM(1) = to_sfixed(-13.2500,QstateIM(1)) then
				char1IM <= "-13.2500";
			elsif QstateIM(1) = to_sfixed(-13.1875,QstateIM(1)) then
				char1IM <= "-13.1875";
			elsif QstateIM(1) = to_sfixed(-13.1250,QstateIM(1)) then
				char1IM <= "-13.1250";
			elsif QstateIM(1) = to_sfixed(-13.0625,QstateIM(1)) then
				char1IM <= "-13.0625";
			elsif QstateIM(1) = to_sfixed(-13.0000,QstateIM(1)) then
				char1IM <= "-13.0000";
			elsif QstateIM(1) = to_sfixed(-12.9375,QstateIM(1)) then
				char1IM <= "-12.9375";
			elsif QstateIM(1) = to_sfixed(-12.8750,QstateIM(1)) then
				char1IM <= "-12.8750";
			elsif QstateIM(1) = to_sfixed(-12.8125,QstateIM(1)) then
				char1IM <= "-12.8125";
			elsif QstateIM(1) = to_sfixed(-12.7500,QstateIM(1)) then
				char1IM <= "-12.7500";
			elsif QstateIM(1) = to_sfixed(-12.6875,QstateIM(1)) then
				char1IM <= "-12.6875";
			elsif QstateIM(1) = to_sfixed(-12.6250,QstateIM(1)) then
				char1IM <= "-12.6250";
			elsif QstateIM(1) = to_sfixed(-12.5625,QstateIM(1)) then
				char1IM <= "-12.5625";
			elsif QstateIM(1) = to_sfixed(-12.5000,QstateIM(1)) then
				char1IM <= "-12.5000";
			elsif QstateIM(1) = to_sfixed(-12.4375,QstateIM(1)) then
				char1IM <= "-12.4375";
			elsif QstateIM(1) = to_sfixed(-12.3750,QstateIM(1)) then
				char1IM <= "-12.3750";
			elsif QstateIM(1) = to_sfixed(-12.3125,QstateIM(1)) then
				char1IM <= "-12.3125";
			elsif QstateIM(1) = to_sfixed(-12.2500,QstateIM(1)) then
				char1IM <= "-12.2500";
			elsif QstateIM(1) = to_sfixed(-12.1875,QstateIM(1)) then
				char1IM <= "-12.1875";
			elsif QstateIM(1) = to_sfixed(-12.1250,QstateIM(1)) then
				char1IM <= "-12.1250";
			elsif QstateIM(1) = to_sfixed(-12.0625,QstateIM(1)) then
				char1IM <= "-12.0625";
			elsif QstateIM(1) = to_sfixed(-12.0000,QstateIM(1)) then
				char1IM <= "-12.0000";
			elsif QstateIM(1) = to_sfixed(-11.9375,QstateIM(1)) then
				char1IM <= "-11.9375";
			elsif QstateIM(1) = to_sfixed(-11.8750,QstateIM(1)) then
				char1IM <= "-11.8750";
			elsif QstateIM(1) = to_sfixed(-11.8125,QstateIM(1)) then
				char1IM <= "-11.8125";
			elsif QstateIM(1) = to_sfixed(-11.7500,QstateIM(1)) then
				char1IM <= "-11.7500";
			elsif QstateIM(1) = to_sfixed(-11.6875,QstateIM(1)) then
				char1IM <= "-11.6875";
			elsif QstateIM(1) = to_sfixed(-11.6250,QstateIM(1)) then
				char1IM <= "-11.6250";
			elsif QstateIM(1) = to_sfixed(-11.5625,QstateIM(1)) then
				char1IM <= "-11.5625";
			elsif QstateIM(1) = to_sfixed(-11.5000,QstateIM(1)) then
				char1IM <= "-11.5000";
			elsif QstateIM(1) = to_sfixed(-11.4375,QstateIM(1)) then
				char1IM <= "-11.4375";
			elsif QstateIM(1) = to_sfixed(-11.3750,QstateIM(1)) then
				char1IM <= "-11.3750";
			elsif QstateIM(1) = to_sfixed(-11.3125,QstateIM(1)) then
				char1IM <= "-11.3125";
			elsif QstateIM(1) = to_sfixed(-11.2500,QstateIM(1)) then
				char1IM <= "-11.2500";
			elsif QstateIM(1) = to_sfixed(-11.1875,QstateIM(1)) then
				char1IM <= "-11.1875";
			elsif QstateIM(1) = to_sfixed(-11.1250,QstateIM(1)) then
				char1IM <= "-11.1250";
			elsif QstateIM(1) = to_sfixed(-11.0625,QstateIM(1)) then
				char1IM <= "-11.0625";
			elsif QstateIM(1) = to_sfixed(-11.0000,QstateIM(1)) then
				char1IM <= "-11.0000";
			elsif QstateIM(1) = to_sfixed(-10.9375,QstateIM(1)) then
				char1IM <= "-10.9375";
			elsif QstateIM(1) = to_sfixed(-10.8750,QstateIM(1)) then
				char1IM <= "-10.8750";
			elsif QstateIM(1) = to_sfixed(-10.8125,QstateIM(1)) then
				char1IM <= "-10.8125";
			elsif QstateIM(1) = to_sfixed(-10.7500,QstateIM(1)) then
				char1IM <= "-10.7500";
			elsif QstateIM(1) = to_sfixed(-10.6875,QstateIM(1)) then
				char1IM <= "-10.6875";
			elsif QstateIM(1) = to_sfixed(-10.6250,QstateIM(1)) then
				char1IM <= "-10.6250";
			elsif QstateIM(1) = to_sfixed(-10.5625,QstateIM(1)) then
				char1IM <= "-10.5625";
			elsif QstateIM(1) = to_sfixed(-10.5000,QstateIM(1)) then
				char1IM <= "-10.5000";
			elsif QstateIM(1) = to_sfixed(-10.4375,QstateIM(1)) then
				char1IM <= "-10.4375";
			elsif QstateIM(1) = to_sfixed(-10.3750,QstateIM(1)) then
				char1IM <= "-10.3750";
			elsif QstateIM(1) = to_sfixed(-10.3125,QstateIM(1)) then
				char1IM <= "-10.3125";
			elsif QstateIM(1) = to_sfixed(-10.2500,QstateIM(1)) then
				char1IM <= "-10.2500";
			elsif QstateIM(1) = to_sfixed(-10.1875,QstateIM(1)) then
				char1IM <= "-10.1875";
			elsif QstateIM(1) = to_sfixed(-10.1250,QstateIM(1)) then
				char1IM <= "-10.1250";
			elsif QstateIM(1) = to_sfixed(-10.0625,QstateIM(1)) then
				char1IM <= "-10.0625";
			elsif QstateIM(1) = to_sfixed(-10.0000,QstateIM(1)) then
				char1IM <= "-10.0000";
			elsif QstateIM(1) = to_sfixed(-9.9375,QstateIM(1)) then
				char1IM <= "--9.9375";
			elsif QstateIM(1) = to_sfixed(-9.8750,QstateIM(1)) then
				char1IM <= "--9.8750";
			elsif QstateIM(1) = to_sfixed(-9.8125,QstateIM(1)) then
				char1IM <= "--9.8125";
			elsif QstateIM(1) = to_sfixed(-9.7500,QstateIM(1)) then
				char1IM <= "--9.7500";
			elsif QstateIM(1) = to_sfixed(-9.6875,QstateIM(1)) then
				char1IM <= "--9.6875";
			elsif QstateIM(1) = to_sfixed(-9.6250,QstateIM(1)) then
				char1IM <= "--9.6250";
			elsif QstateIM(1) = to_sfixed(-9.5625,QstateIM(1)) then
				char1IM <= "--9.5625";
			elsif QstateIM(1) = to_sfixed(-9.5000,QstateIM(1)) then
				char1IM <= "--9.5000";
			elsif QstateIM(1) = to_sfixed(-9.4375,QstateIM(1)) then
				char1IM <= "--9.4375";
			elsif QstateIM(1) = to_sfixed(-9.3750,QstateIM(1)) then
				char1IM <= "--9.3750";
			elsif QstateIM(1) = to_sfixed(-9.3125,QstateIM(1)) then
				char1IM <= "--9.3125";
			elsif QstateIM(1) = to_sfixed(-9.2500,QstateIM(1)) then
				char1IM <= "--9.2500";
			elsif QstateIM(1) = to_sfixed(-9.1875,QstateIM(1)) then
				char1IM <= "--9.1875";
			elsif QstateIM(1) = to_sfixed(-9.1250,QstateIM(1)) then
				char1IM <= "--9.1250";
			elsif QstateIM(1) = to_sfixed(-9.0625,QstateIM(1)) then
				char1IM <= "--9.0625";
			elsif QstateIM(1) = to_sfixed(-9.0000,QstateIM(1)) then
				char1IM <= "--9.0000";
			elsif QstateIM(1) = to_sfixed(-8.9375,QstateIM(1)) then
				char1IM <= "--8.9375";
			elsif QstateIM(1) = to_sfixed(-8.8750,QstateIM(1)) then
				char1IM <= "--8.8750";
			elsif QstateIM(1) = to_sfixed(-8.8125,QstateIM(1)) then
				char1IM <= "--8.8125";
			elsif QstateIM(1) = to_sfixed(-8.7500,QstateIM(1)) then
				char1IM <= "--8.7500";
			elsif QstateIM(1) = to_sfixed(-8.6875,QstateIM(1)) then
				char1IM <= "--8.6875";
			elsif QstateIM(1) = to_sfixed(-8.6250,QstateIM(1)) then
				char1IM <= "--8.6250";
			elsif QstateIM(1) = to_sfixed(-8.5625,QstateIM(1)) then
				char1IM <= "--8.5625";
			elsif QstateIM(1) = to_sfixed(-8.5000,QstateIM(1)) then
				char1IM <= "--8.5000";
			elsif QstateIM(1) = to_sfixed(-8.4375,QstateIM(1)) then
				char1IM <= "--8.4375";
			elsif QstateIM(1) = to_sfixed(-8.3750,QstateIM(1)) then
				char1IM <= "--8.3750";
			elsif QstateIM(1) = to_sfixed(-8.3125,QstateIM(1)) then
				char1IM <= "--8.3125";
			elsif QstateIM(1) = to_sfixed(-8.2500,QstateIM(1)) then
				char1IM <= "--8.2500";
			elsif QstateIM(1) = to_sfixed(-8.1875,QstateIM(1)) then
				char1IM <= "--8.1875";
			elsif QstateIM(1) = to_sfixed(-8.1250,QstateIM(1)) then
				char1IM <= "--8.1250";
			elsif QstateIM(1) = to_sfixed(-8.0625,QstateIM(1)) then
				char1IM <= "--8.0625";
			elsif QstateIM(1) = to_sfixed(-8.0000,QstateIM(1)) then
				char1IM <= "--8.0000";
			elsif QstateIM(1) = to_sfixed(-7.9375,QstateIM(1)) then
				char1IM <= "--7.9375";
			elsif QstateIM(1) = to_sfixed(-7.8750,QstateIM(1)) then
				char1IM <= "--7.8750";
			elsif QstateIM(1) = to_sfixed(-7.8125,QstateIM(1)) then
				char1IM <= "--7.8125";
			elsif QstateIM(1) = to_sfixed(-7.7500,QstateIM(1)) then
				char1IM <= "--7.7500";
			elsif QstateIM(1) = to_sfixed(-7.6875,QstateIM(1)) then
				char1IM <= "--7.6875";
			elsif QstateIM(1) = to_sfixed(-7.6250,QstateIM(1)) then
				char1IM <= "--7.6250";
			elsif QstateIM(1) = to_sfixed(-7.5625,QstateIM(1)) then
				char1IM <= "--7.5625";
			elsif QstateIM(1) = to_sfixed(-7.5000,QstateIM(1)) then
				char1IM <= "--7.5000";
			elsif QstateIM(1) = to_sfixed(-7.4375,QstateIM(1)) then
				char1IM <= "--7.4375";
			elsif QstateIM(1) = to_sfixed(-7.3750,QstateIM(1)) then
				char1IM <= "--7.3750";
			elsif QstateIM(1) = to_sfixed(-7.3125,QstateIM(1)) then
				char1IM <= "--7.3125";
			elsif QstateIM(1) = to_sfixed(-7.2500,QstateIM(1)) then
				char1IM <= "--7.2500";
			elsif QstateIM(1) = to_sfixed(-7.1875,QstateIM(1)) then
				char1IM <= "--7.1875";
			elsif QstateIM(1) = to_sfixed(-7.1250,QstateIM(1)) then
				char1IM <= "--7.1250";
			elsif QstateIM(1) = to_sfixed(-7.0625,QstateIM(1)) then
				char1IM <= "--7.0625";
			elsif QstateIM(1) = to_sfixed(-7.0000,QstateIM(1)) then
				char1IM <= "--7.0000";
			elsif QstateIM(1) = to_sfixed(-6.9375,QstateIM(1)) then
				char1IM <= "--6.9375";
			elsif QstateIM(1) = to_sfixed(-6.8750,QstateIM(1)) then
				char1IM <= "--6.8750";
			elsif QstateIM(1) = to_sfixed(-6.8125,QstateIM(1)) then
				char1IM <= "--6.8125";
			elsif QstateIM(1) = to_sfixed(-6.7500,QstateIM(1)) then
				char1IM <= "--6.7500";
			elsif QstateIM(1) = to_sfixed(-6.6875,QstateIM(1)) then
				char1IM <= "--6.6875";
			elsif QstateIM(1) = to_sfixed(-6.6250,QstateIM(1)) then
				char1IM <= "--6.6250";
			elsif QstateIM(1) = to_sfixed(-6.5625,QstateIM(1)) then
				char1IM <= "--6.5625";
			elsif QstateIM(1) = to_sfixed(-6.5000,QstateIM(1)) then
				char1IM <= "--6.5000";
			elsif QstateIM(1) = to_sfixed(-6.4375,QstateIM(1)) then
				char1IM <= "--6.4375";
			elsif QstateIM(1) = to_sfixed(-6.3750,QstateIM(1)) then
				char1IM <= "--6.3750";
			elsif QstateIM(1) = to_sfixed(-6.3125,QstateIM(1)) then
				char1IM <= "--6.3125";
			elsif QstateIM(1) = to_sfixed(-6.2500,QstateIM(1)) then
				char1IM <= "--6.2500";
			elsif QstateIM(1) = to_sfixed(-6.1875,QstateIM(1)) then
				char1IM <= "--6.1875";
			elsif QstateIM(1) = to_sfixed(-6.1250,QstateIM(1)) then
				char1IM <= "--6.1250";
			elsif QstateIM(1) = to_sfixed(-6.0625,QstateIM(1)) then
				char1IM <= "--6.0625";
			elsif QstateIM(1) = to_sfixed(-6.0000,QstateIM(1)) then
				char1IM <= "--6.0000";
			elsif QstateIM(1) = to_sfixed(-5.9375,QstateIM(1)) then
				char1IM <= "--5.9375";
			elsif QstateIM(1) = to_sfixed(-5.8750,QstateIM(1)) then
				char1IM <= "--5.8750";
			elsif QstateIM(1) = to_sfixed(-5.8125,QstateIM(1)) then
				char1IM <= "--5.8125";
			elsif QstateIM(1) = to_sfixed(-5.7500,QstateIM(1)) then
				char1IM <= "--5.7500";
			elsif QstateIM(1) = to_sfixed(-5.6875,QstateIM(1)) then
				char1IM <= "--5.6875";
			elsif QstateIM(1) = to_sfixed(-5.6250,QstateIM(1)) then
				char1IM <= "--5.6250";
			elsif QstateIM(1) = to_sfixed(-5.5625,QstateIM(1)) then
				char1IM <= "--5.5625";
			elsif QstateIM(1) = to_sfixed(-5.5000,QstateIM(1)) then
				char1IM <= "--5.5000";
			elsif QstateIM(1) = to_sfixed(-5.4375,QstateIM(1)) then
				char1IM <= "--5.4375";
			elsif QstateIM(1) = to_sfixed(-5.3750,QstateIM(1)) then
				char1IM <= "--5.3750";
			elsif QstateIM(1) = to_sfixed(-5.3125,QstateIM(1)) then
				char1IM <= "--5.3125";
			elsif QstateIM(1) = to_sfixed(-5.2500,QstateIM(1)) then
				char1IM <= "--5.2500";
			elsif QstateIM(1) = to_sfixed(-5.1875,QstateIM(1)) then
				char1IM <= "--5.1875";
			elsif QstateIM(1) = to_sfixed(-5.1250,QstateIM(1)) then
				char1IM <= "--5.1250";
			elsif QstateIM(1) = to_sfixed(-5.0625,QstateIM(1)) then
				char1IM <= "--5.0625";
			elsif QstateIM(1) = to_sfixed(-5.0000,QstateIM(1)) then
				char1IM <= "--5.0000";
			elsif QstateIM(1) = to_sfixed(-4.9375,QstateIM(1)) then
				char1IM <= "--4.9375";
			elsif QstateIM(1) = to_sfixed(-4.8750,QstateIM(1)) then
				char1IM <= "--4.8750";
			elsif QstateIM(1) = to_sfixed(-4.8125,QstateIM(1)) then
				char1IM <= "--4.8125";
			elsif QstateIM(1) = to_sfixed(-4.7500,QstateIM(1)) then
				char1IM <= "--4.7500";
			elsif QstateIM(1) = to_sfixed(-4.6875,QstateIM(1)) then
				char1IM <= "--4.6875";
			elsif QstateIM(1) = to_sfixed(-4.6250,QstateIM(1)) then
				char1IM <= "--4.6250";
			elsif QstateIM(1) = to_sfixed(-4.5625,QstateIM(1)) then
				char1IM <= "--4.5625";
			elsif QstateIM(1) = to_sfixed(-4.5000,QstateIM(1)) then
				char1IM <= "--4.5000";
			elsif QstateIM(1) = to_sfixed(-4.4375,QstateIM(1)) then
				char1IM <= "--4.4375";
			elsif QstateIM(1) = to_sfixed(-4.3750,QstateIM(1)) then
				char1IM <= "--4.3750";
			elsif QstateIM(1) = to_sfixed(-4.3125,QstateIM(1)) then
				char1IM <= "--4.3125";
			elsif QstateIM(1) = to_sfixed(-4.2500,QstateIM(1)) then
				char1IM <= "--4.2500";
			elsif QstateIM(1) = to_sfixed(-4.1875,QstateIM(1)) then
				char1IM <= "--4.1875";
			elsif QstateIM(1) = to_sfixed(-4.1250,QstateIM(1)) then
				char1IM <= "--4.1250";
			elsif QstateIM(1) = to_sfixed(-4.0625,QstateIM(1)) then
				char1IM <= "--4.0625";
			elsif QstateIM(1) = to_sfixed(-4.0000,QstateIM(1)) then
				char1IM <= "--4.0000";
			elsif QstateIM(1) = to_sfixed(-3.9375,QstateIM(1)) then
				char1IM <= "--3.9375";
			elsif QstateIM(1) = to_sfixed(-3.8750,QstateIM(1)) then
				char1IM <= "--3.8750";
			elsif QstateIM(1) = to_sfixed(-3.8125,QstateIM(1)) then
				char1IM <= "--3.8125";
			elsif QstateIM(1) = to_sfixed(-3.7500,QstateIM(1)) then
				char1IM <= "--3.7500";
			elsif QstateIM(1) = to_sfixed(-3.6875,QstateIM(1)) then
				char1IM <= "--3.6875";
			elsif QstateIM(1) = to_sfixed(-3.6250,QstateIM(1)) then
				char1IM <= "--3.6250";
			elsif QstateIM(1) = to_sfixed(-3.5625,QstateIM(1)) then
				char1IM <= "--3.5625";
			elsif QstateIM(1) = to_sfixed(-3.5000,QstateIM(1)) then
				char1IM <= "--3.5000";
			elsif QstateIM(1) = to_sfixed(-3.4375,QstateIM(1)) then
				char1IM <= "--3.4375";
			elsif QstateIM(1) = to_sfixed(-3.3750,QstateIM(1)) then
				char1IM <= "--3.3750";
			elsif QstateIM(1) = to_sfixed(-3.3125,QstateIM(1)) then
				char1IM <= "--3.3125";
			elsif QstateIM(1) = to_sfixed(-3.2500,QstateIM(1)) then
				char1IM <= "--3.2500";
			elsif QstateIM(1) = to_sfixed(-3.1875,QstateIM(1)) then
				char1IM <= "--3.1875";
			elsif QstateIM(1) = to_sfixed(-3.1250,QstateIM(1)) then
				char1IM <= "--3.1250";
			elsif QstateIM(1) = to_sfixed(-3.0625,QstateIM(1)) then
				char1IM <= "--3.0625";
			elsif QstateIM(1) = to_sfixed(-3.0000,QstateIM(1)) then
				char1IM <= "--3.0000";
			elsif QstateIM(1) = to_sfixed(-2.9375,QstateIM(1)) then
				char1IM <= "--2.9375";
			elsif QstateIM(1) = to_sfixed(-2.8750,QstateIM(1)) then
				char1IM <= "--2.8750";
			elsif QstateIM(1) = to_sfixed(-2.8125,QstateIM(1)) then
				char1IM <= "--2.8125";
			elsif QstateIM(1) = to_sfixed(-2.7500,QstateIM(1)) then
				char1IM <= "--2.7500";
			elsif QstateIM(1) = to_sfixed(-2.6875,QstateIM(1)) then
				char1IM <= "--2.6875";
			elsif QstateIM(1) = to_sfixed(-2.6250,QstateIM(1)) then
				char1IM <= "--2.6250";
			elsif QstateIM(1) = to_sfixed(-2.5625,QstateIM(1)) then
				char1IM <= "--2.5625";
			elsif QstateIM(1) = to_sfixed(-2.5000,QstateIM(1)) then
				char1IM <= "--2.5000";
			elsif QstateIM(1) = to_sfixed(-2.4375,QstateIM(1)) then
				char1IM <= "--2.4375";
			elsif QstateIM(1) = to_sfixed(-2.3750,QstateIM(1)) then
				char1IM <= "--2.3750";
			elsif QstateIM(1) = to_sfixed(-2.3125,QstateIM(1)) then
				char1IM <= "--2.3125";
			elsif QstateIM(1) = to_sfixed(-2.2500,QstateIM(1)) then
				char1IM <= "--2.2500";
			elsif QstateIM(1) = to_sfixed(-2.1875,QstateIM(1)) then
				char1IM <= "--2.1875";
			elsif QstateIM(1) = to_sfixed(-2.1250,QstateIM(1)) then
				char1IM <= "--2.1250";
			elsif QstateIM(1) = to_sfixed(-2.0625,QstateIM(1)) then
				char1IM <= "--2.0625";
			elsif QstateIM(1) = to_sfixed(-2.0000,QstateIM(1)) then
				char1IM <= "--2.0000";
			elsif QstateIM(1) = to_sfixed(-1.9375,QstateIM(1)) then
				char1IM <= "--1.9375";
			elsif QstateIM(1) = to_sfixed(-1.8750,QstateIM(1)) then
				char1IM <= "--1.8750";
			elsif QstateIM(1) = to_sfixed(-1.8125,QstateIM(1)) then
				char1IM <= "--1.8125";
			elsif QstateIM(1) = to_sfixed(-1.7500,QstateIM(1)) then
				char1IM <= "--1.7500";
			elsif QstateIM(1) = to_sfixed(-1.6875,QstateIM(1)) then
				char1IM <= "--1.6875";
			elsif QstateIM(1) = to_sfixed(-1.6250,QstateIM(1)) then
				char1IM <= "--1.6250";
			elsif QstateIM(1) = to_sfixed(-1.5625,QstateIM(1)) then
				char1IM <= "--1.5625";
			elsif QstateIM(1) = to_sfixed(-1.5000,QstateIM(1)) then
				char1IM <= "--1.5000";
			elsif QstateIM(1) = to_sfixed(-1.4375,QstateIM(1)) then
				char1IM <= "--1.4375";
			elsif QstateIM(1) = to_sfixed(-1.3750,QstateIM(1)) then
				char1IM <= "--1.3750";
			elsif QstateIM(1) = to_sfixed(-1.3125,QstateIM(1)) then
				char1IM <= "--1.3125";
			elsif QstateIM(1) = to_sfixed(-1.2500,QstateIM(1)) then
				char1IM <= "--1.2500";
			elsif QstateIM(1) = to_sfixed(-1.1875,QstateIM(1)) then
				char1IM <= "--1.1875";
			elsif QstateIM(1) = to_sfixed(-1.1250,QstateIM(1)) then
				char1IM <= "--1.1250";
			elsif QstateIM(1) = to_sfixed(-1.0625,QstateIM(1)) then
				char1IM <= "--1.0625";
			elsif QstateIM(1) = to_sfixed(-1.0000,QstateIM(1)) then
				char1IM <= "--1.0000";
			elsif QstateIM(1) = to_sfixed(-0.9375,QstateIM(1)) then
				char1IM <= "--0.9375";
			elsif QstateIM(1) = to_sfixed(-0.8750,QstateIM(1)) then
				char1IM <= "--0.8750";
			elsif QstateIM(1) = to_sfixed(-0.8125,QstateIM(1)) then
				char1IM <= "--0.8125";
			elsif QstateIM(1) = to_sfixed(-0.7500,QstateIM(1)) then
				char1IM <= "--0.7500";
			elsif QstateIM(1) = to_sfixed(-0.6875,QstateIM(1)) then
				char1IM <= "--0.6875";
			elsif QstateIM(1) = to_sfixed(-0.6250,QstateIM(1)) then
				char1IM <= "--0.6250";
			elsif QstateIM(1) = to_sfixed(-0.5625,QstateIM(1)) then
				char1IM <= "--0.5625";
			elsif QstateIM(1) = to_sfixed(-0.5000,QstateIM(1)) then
				char1IM <= "--0.5000";
			elsif QstateIM(1) = to_sfixed(-0.4375,QstateIM(1)) then
				char1IM <= "--0.4375";
			elsif QstateIM(1) = to_sfixed(-0.3750,QstateIM(1)) then
				char1IM <= "--0.3750";
			elsif QstateIM(1) = to_sfixed(-0.3125,QstateIM(1)) then
				char1IM <= "--0.3125";
			elsif QstateIM(1) = to_sfixed(-0.2500,QstateIM(1)) then
				char1IM <= "--0.2500";
			elsif QstateIM(1) = to_sfixed(-0.1875,QstateIM(1)) then
				char1IM <= "--0.1875";
			elsif QstateIM(1) = to_sfixed(-0.1250,QstateIM(1)) then
				char1IM <= "--0.1250";
			elsif QstateIM(1) = to_sfixed(-0.0625,QstateIM(1)) then
				char1IM <= "--0.0625";
			elsif QstateIM(1) = to_sfixed(00.0000,QstateIM(1)) then
				char1IM <= "+00.0000";
			elsif QstateIM(1) = to_sfixed(00.0625,QstateIM(1)) then
				char1IM <= "+00.0625";
			elsif QstateIM(1) = to_sfixed(00.1250,QstateIM(1)) then
				char1IM <= "+00.1250";
			elsif QstateIM(1) = to_sfixed(00.1875,QstateIM(1)) then
				char1IM <= "+00.1875";
			elsif QstateIM(1) = to_sfixed(00.2500,QstateIM(1)) then
				char1IM <= "+00.2500";
			elsif QstateIM(1) = to_sfixed(00.3125,QstateIM(1)) then
				char1IM <= "+00.3125";
			elsif QstateIM(1) = to_sfixed(00.3750,QstateIM(1)) then
				char1IM <= "+00.3750";
			elsif QstateIM(1) = to_sfixed(00.4375,QstateIM(1)) then
				char1IM <= "+00.4375";
			elsif QstateIM(1) = to_sfixed(00.5000,QstateIM(1)) then
				char1IM <= "+00.5000";
			elsif QstateIM(1) = to_sfixed(00.5625,QstateIM(1)) then
				char1IM <= "+00.5625";
			elsif QstateIM(1) = to_sfixed(00.6250,QstateIM(1)) then
				char1IM <= "+00.6250";
			elsif QstateIM(1) = to_sfixed(00.6875,QstateIM(1)) then
				char1IM <= "+00.6875";
			elsif QstateIM(1) = to_sfixed(00.7500,QstateIM(1)) then
				char1IM <= "+00.7500";
			elsif QstateIM(1) = to_sfixed(00.8125,QstateIM(1)) then
				char1IM <= "+00.8125";
			elsif QstateIM(1) = to_sfixed(00.8750,QstateIM(1)) then
				char1IM <= "+00.8750";
			elsif QstateIM(1) = to_sfixed(00.9375,QstateIM(1)) then
				char1IM <= "+00.9375";
			elsif QstateIM(1) = to_sfixed(01.0000,QstateIM(1)) then
				char1IM <= "+01.0000";
			elsif QstateIM(1) = to_sfixed(01.0625,QstateIM(1)) then
				char1IM <= "+01.0625";
			elsif QstateIM(1) = to_sfixed(01.1250,QstateIM(1)) then
				char1IM <= "+01.1250";
			elsif QstateIM(1) = to_sfixed(01.1875,QstateIM(1)) then
				char1IM <= "+01.1875";
			elsif QstateIM(1) = to_sfixed(01.2500,QstateIM(1)) then
				char1IM <= "+01.2500";
			elsif QstateIM(1) = to_sfixed(01.3125,QstateIM(1)) then
				char1IM <= "+01.3125";
			elsif QstateIM(1) = to_sfixed(01.3750,QstateIM(1)) then
				char1IM <= "+01.3750";
			elsif QstateIM(1) = to_sfixed(01.4375,QstateIM(1)) then
				char1IM <= "+01.4375";
			elsif QstateIM(1) = to_sfixed(01.5000,QstateIM(1)) then
				char1IM <= "+01.5000";
			elsif QstateIM(1) = to_sfixed(01.5625,QstateIM(1)) then
				char1IM <= "+01.5625";
			elsif QstateIM(1) = to_sfixed(01.6250,QstateIM(1)) then
				char1IM <= "+01.6250";
			elsif QstateIM(1) = to_sfixed(01.6875,QstateIM(1)) then
				char1IM <= "+01.6875";
			elsif QstateIM(1) = to_sfixed(01.7500,QstateIM(1)) then
				char1IM <= "+01.7500";
			elsif QstateIM(1) = to_sfixed(01.8125,QstateIM(1)) then
				char1IM <= "+01.8125";
			elsif QstateIM(1) = to_sfixed(01.8750,QstateIM(1)) then
				char1IM <= "+01.8750";
			elsif QstateIM(1) = to_sfixed(01.9375,QstateIM(1)) then
				char1IM <= "+01.9375";
			elsif QstateIM(1) = to_sfixed(02.0000,QstateIM(1)) then
				char1IM <= "+02.0000";
			elsif QstateIM(1) = to_sfixed(02.0625,QstateIM(1)) then
				char1IM <= "+02.0625";
			elsif QstateIM(1) = to_sfixed(02.1250,QstateIM(1)) then
				char1IM <= "+02.1250";
			elsif QstateIM(1) = to_sfixed(02.1875,QstateIM(1)) then
				char1IM <= "+02.1875";
			elsif QstateIM(1) = to_sfixed(02.2500,QstateIM(1)) then
				char1IM <= "+02.2500";
			elsif QstateIM(1) = to_sfixed(02.3125,QstateIM(1)) then
				char1IM <= "+02.3125";
			elsif QstateIM(1) = to_sfixed(02.3750,QstateIM(1)) then
				char1IM <= "+02.3750";
			elsif QstateIM(1) = to_sfixed(02.4375,QstateIM(1)) then
				char1IM <= "+02.4375";
			elsif QstateIM(1) = to_sfixed(02.5000,QstateIM(1)) then
				char1IM <= "+02.5000";
			elsif QstateIM(1) = to_sfixed(02.5625,QstateIM(1)) then
				char1IM <= "+02.5625";
			elsif QstateIM(1) = to_sfixed(02.6250,QstateIM(1)) then
				char1IM <= "+02.6250";
			elsif QstateIM(1) = to_sfixed(02.6875,QstateIM(1)) then
				char1IM <= "+02.6875";
			elsif QstateIM(1) = to_sfixed(02.7500,QstateIM(1)) then
				char1IM <= "+02.7500";
			elsif QstateIM(1) = to_sfixed(02.8125,QstateIM(1)) then
				char1IM <= "+02.8125";
			elsif QstateIM(1) = to_sfixed(02.8750,QstateIM(1)) then
				char1IM <= "+02.8750";
			elsif QstateIM(1) = to_sfixed(02.9375,QstateIM(1)) then
				char1IM <= "+02.9375";
			elsif QstateIM(1) = to_sfixed(03.0000,QstateIM(1)) then
				char1IM <= "+03.0000";
			elsif QstateIM(1) = to_sfixed(03.0625,QstateIM(1)) then
				char1IM <= "+03.0625";
			elsif QstateIM(1) = to_sfixed(03.1250,QstateIM(1)) then
				char1IM <= "+03.1250";
			elsif QstateIM(1) = to_sfixed(03.1875,QstateIM(1)) then
				char1IM <= "+03.1875";
			elsif QstateIM(1) = to_sfixed(03.2500,QstateIM(1)) then
				char1IM <= "+03.2500";
			elsif QstateIM(1) = to_sfixed(03.3125,QstateIM(1)) then
				char1IM <= "+03.3125";
			elsif QstateIM(1) = to_sfixed(03.3750,QstateIM(1)) then
				char1IM <= "+03.3750";
			elsif QstateIM(1) = to_sfixed(03.4375,QstateIM(1)) then
				char1IM <= "+03.4375";
			elsif QstateIM(1) = to_sfixed(03.5000,QstateIM(1)) then
				char1IM <= "+03.5000";
			elsif QstateIM(1) = to_sfixed(03.5625,QstateIM(1)) then
				char1IM <= "+03.5625";
			elsif QstateIM(1) = to_sfixed(03.6250,QstateIM(1)) then
				char1IM <= "+03.6250";
			elsif QstateIM(1) = to_sfixed(03.6875,QstateIM(1)) then
				char1IM <= "+03.6875";
			elsif QstateIM(1) = to_sfixed(03.7500,QstateIM(1)) then
				char1IM <= "+03.7500";
			elsif QstateIM(1) = to_sfixed(03.8125,QstateIM(1)) then
				char1IM <= "+03.8125";
			elsif QstateIM(1) = to_sfixed(03.8750,QstateIM(1)) then
				char1IM <= "+03.8750";
			elsif QstateIM(1) = to_sfixed(03.9375,QstateIM(1)) then
				char1IM <= "+03.9375";
			elsif QstateIM(1) = to_sfixed(04.0000,QstateIM(1)) then
				char1IM <= "+04.0000";
			elsif QstateIM(1) = to_sfixed(04.0625,QstateIM(1)) then
				char1IM <= "+04.0625";
			elsif QstateIM(1) = to_sfixed(04.1250,QstateIM(1)) then
				char1IM <= "+04.1250";
			elsif QstateIM(1) = to_sfixed(04.1875,QstateIM(1)) then
				char1IM <= "+04.1875";
			elsif QstateIM(1) = to_sfixed(04.2500,QstateIM(1)) then
				char1IM <= "+04.2500";
			elsif QstateIM(1) = to_sfixed(04.3125,QstateIM(1)) then
				char1IM <= "+04.3125";
			elsif QstateIM(1) = to_sfixed(04.3750,QstateIM(1)) then
				char1IM <= "+04.3750";
			elsif QstateIM(1) = to_sfixed(04.4375,QstateIM(1)) then
				char1IM <= "+04.4375";
			elsif QstateIM(1) = to_sfixed(04.5000,QstateIM(1)) then
				char1IM <= "+04.5000";
			elsif QstateIM(1) = to_sfixed(04.5625,QstateIM(1)) then
				char1IM <= "+04.5625";
			elsif QstateIM(1) = to_sfixed(04.6250,QstateIM(1)) then
				char1IM <= "+04.6250";
			elsif QstateIM(1) = to_sfixed(04.6875,QstateIM(1)) then
				char1IM <= "+04.6875";
			elsif QstateIM(1) = to_sfixed(04.7500,QstateIM(1)) then
				char1IM <= "+04.7500";
			elsif QstateIM(1) = to_sfixed(04.8125,QstateIM(1)) then
				char1IM <= "+04.8125";
			elsif QstateIM(1) = to_sfixed(04.8750,QstateIM(1)) then
				char1IM <= "+04.8750";
			elsif QstateIM(1) = to_sfixed(04.9375,QstateIM(1)) then
				char1IM <= "+04.9375";
			elsif QstateIM(1) = to_sfixed(05.0000,QstateIM(1)) then
				char1IM <= "+05.0000";
			elsif QstateIM(1) = to_sfixed(05.0625,QstateIM(1)) then
				char1IM <= "+05.0625";
			elsif QstateIM(1) = to_sfixed(05.1250,QstateIM(1)) then
				char1IM <= "+05.1250";
			elsif QstateIM(1) = to_sfixed(05.1875,QstateIM(1)) then
				char1IM <= "+05.1875";
			elsif QstateIM(1) = to_sfixed(05.2500,QstateIM(1)) then
				char1IM <= "+05.2500";
			elsif QstateIM(1) = to_sfixed(05.3125,QstateIM(1)) then
				char1IM <= "+05.3125";
			elsif QstateIM(1) = to_sfixed(05.3750,QstateIM(1)) then
				char1IM <= "+05.3750";
			elsif QstateIM(1) = to_sfixed(05.4375,QstateIM(1)) then
				char1IM <= "+05.4375";
			elsif QstateIM(1) = to_sfixed(05.5000,QstateIM(1)) then
				char1IM <= "+05.5000";
			elsif QstateIM(1) = to_sfixed(05.5625,QstateIM(1)) then
				char1IM <= "+05.5625";
			elsif QstateIM(1) = to_sfixed(05.6250,QstateIM(1)) then
				char1IM <= "+05.6250";
			elsif QstateIM(1) = to_sfixed(05.6875,QstateIM(1)) then
				char1IM <= "+05.6875";
			elsif QstateIM(1) = to_sfixed(05.7500,QstateIM(1)) then
				char1IM <= "+05.7500";
			elsif QstateIM(1) = to_sfixed(05.8125,QstateIM(1)) then
				char1IM <= "+05.8125";
			elsif QstateIM(1) = to_sfixed(05.8750,QstateIM(1)) then
				char1IM <= "+05.8750";
			elsif QstateIM(1) = to_sfixed(05.9375,QstateIM(1)) then
				char1IM <= "+05.9375";
			elsif QstateIM(1) = to_sfixed(06.0000,QstateIM(1)) then
				char1IM <= "+06.0000";
			elsif QstateIM(1) = to_sfixed(06.0625,QstateIM(1)) then
				char1IM <= "+06.0625";
			elsif QstateIM(1) = to_sfixed(06.1250,QstateIM(1)) then
				char1IM <= "+06.1250";
			elsif QstateIM(1) = to_sfixed(06.1875,QstateIM(1)) then
				char1IM <= "+06.1875";
			elsif QstateIM(1) = to_sfixed(06.2500,QstateIM(1)) then
				char1IM <= "+06.2500";
			elsif QstateIM(1) = to_sfixed(06.3125,QstateIM(1)) then
				char1IM <= "+06.3125";
			elsif QstateIM(1) = to_sfixed(06.3750,QstateIM(1)) then
				char1IM <= "+06.3750";
			elsif QstateIM(1) = to_sfixed(06.4375,QstateIM(1)) then
				char1IM <= "+06.4375";
			elsif QstateIM(1) = to_sfixed(06.5000,QstateIM(1)) then
				char1IM <= "+06.5000";
			elsif QstateIM(1) = to_sfixed(06.5625,QstateIM(1)) then
				char1IM <= "+06.5625";
			elsif QstateIM(1) = to_sfixed(06.6250,QstateIM(1)) then
				char1IM <= "+06.6250";
			elsif QstateIM(1) = to_sfixed(06.6875,QstateIM(1)) then
				char1IM <= "+06.6875";
			elsif QstateIM(1) = to_sfixed(06.7500,QstateIM(1)) then
				char1IM <= "+06.7500";
			elsif QstateIM(1) = to_sfixed(06.8125,QstateIM(1)) then
				char1IM <= "+06.8125";
			elsif QstateIM(1) = to_sfixed(06.8750,QstateIM(1)) then
				char1IM <= "+06.8750";
			elsif QstateIM(1) = to_sfixed(06.9375,QstateIM(1)) then
				char1IM <= "+06.9375";
			elsif QstateIM(1) = to_sfixed(07.0000,QstateIM(1)) then
				char1IM <= "+07.0000";
			elsif QstateIM(1) = to_sfixed(07.0625,QstateIM(1)) then
				char1IM <= "+07.0625";
			elsif QstateIM(1) = to_sfixed(07.1250,QstateIM(1)) then
				char1IM <= "+07.1250";
			elsif QstateIM(1) = to_sfixed(07.1875,QstateIM(1)) then
				char1IM <= "+07.1875";
			elsif QstateIM(1) = to_sfixed(07.2500,QstateIM(1)) then
				char1IM <= "+07.2500";
			elsif QstateIM(1) = to_sfixed(07.3125,QstateIM(1)) then
				char1IM <= "+07.3125";
			elsif QstateIM(1) = to_sfixed(07.3750,QstateIM(1)) then
				char1IM <= "+07.3750";
			elsif QstateIM(1) = to_sfixed(07.4375,QstateIM(1)) then
				char1IM <= "+07.4375";
			elsif QstateIM(1) = to_sfixed(07.5000,QstateIM(1)) then
				char1IM <= "+07.5000";
			elsif QstateIM(1) = to_sfixed(07.5625,QstateIM(1)) then
				char1IM <= "+07.5625";
			elsif QstateIM(1) = to_sfixed(07.6250,QstateIM(1)) then
				char1IM <= "+07.6250";
			elsif QstateIM(1) = to_sfixed(07.6875,QstateIM(1)) then
				char1IM <= "+07.6875";
			elsif QstateIM(1) = to_sfixed(07.7500,QstateIM(1)) then
				char1IM <= "+07.7500";
			elsif QstateIM(1) = to_sfixed(07.8125,QstateIM(1)) then
				char1IM <= "+07.8125";
			elsif QstateIM(1) = to_sfixed(07.8750,QstateIM(1)) then
				char1IM <= "+07.8750";
			elsif QstateIM(1) = to_sfixed(07.9375,QstateIM(1)) then
				char1IM <= "+07.9375";
			elsif QstateIM(1) = to_sfixed(08.0000,QstateIM(1)) then
				char1IM <= "+08.0000";
			elsif QstateIM(1) = to_sfixed(08.0625,QstateIM(1)) then
				char1IM <= "+08.0625";
			elsif QstateIM(1) = to_sfixed(08.1250,QstateIM(1)) then
				char1IM <= "+08.1250";
			elsif QstateIM(1) = to_sfixed(08.1875,QstateIM(1)) then
				char1IM <= "+08.1875";
			elsif QstateIM(1) = to_sfixed(08.2500,QstateIM(1)) then
				char1IM <= "+08.2500";
			elsif QstateIM(1) = to_sfixed(08.3125,QstateIM(1)) then
				char1IM <= "+08.3125";
			elsif QstateIM(1) = to_sfixed(08.3750,QstateIM(1)) then
				char1IM <= "+08.3750";
			elsif QstateIM(1) = to_sfixed(08.4375,QstateIM(1)) then
				char1IM <= "+08.4375";
			elsif QstateIM(1) = to_sfixed(08.5000,QstateIM(1)) then
				char1IM <= "+08.5000";
			elsif QstateIM(1) = to_sfixed(08.5625,QstateIM(1)) then
				char1IM <= "+08.5625";
			elsif QstateIM(1) = to_sfixed(08.6250,QstateIM(1)) then
				char1IM <= "+08.6250";
			elsif QstateIM(1) = to_sfixed(08.6875,QstateIM(1)) then
				char1IM <= "+08.6875";
			elsif QstateIM(1) = to_sfixed(08.7500,QstateIM(1)) then
				char1IM <= "+08.7500";
			elsif QstateIM(1) = to_sfixed(08.8125,QstateIM(1)) then
				char1IM <= "+08.8125";
			elsif QstateIM(1) = to_sfixed(08.8750,QstateIM(1)) then
				char1IM <= "+08.8750";
			elsif QstateIM(1) = to_sfixed(08.9375,QstateIM(1)) then
				char1IM <= "+08.9375";
			elsif QstateIM(1) = to_sfixed(09.0000,QstateIM(1)) then
				char1IM <= "+09.0000";
			elsif QstateIM(1) = to_sfixed(09.0625,QstateIM(1)) then
				char1IM <= "+09.0625";
			elsif QstateIM(1) = to_sfixed(09.1250,QstateIM(1)) then
				char1IM <= "+09.1250";
			elsif QstateIM(1) = to_sfixed(09.1875,QstateIM(1)) then
				char1IM <= "+09.1875";
			elsif QstateIM(1) = to_sfixed(09.2500,QstateIM(1)) then
				char1IM <= "+09.2500";
			elsif QstateIM(1) = to_sfixed(09.3125,QstateIM(1)) then
				char1IM <= "+09.3125";
			elsif QstateIM(1) = to_sfixed(09.3750,QstateIM(1)) then
				char1IM <= "+09.3750";
			elsif QstateIM(1) = to_sfixed(09.4375,QstateIM(1)) then
				char1IM <= "+09.4375";
			elsif QstateIM(1) = to_sfixed(09.5000,QstateIM(1)) then
				char1IM <= "+09.5000";
			elsif QstateIM(1) = to_sfixed(09.5625,QstateIM(1)) then
				char1IM <= "+09.5625";
			elsif QstateIM(1) = to_sfixed(09.6250,QstateIM(1)) then
				char1IM <= "+09.6250";
			elsif QstateIM(1) = to_sfixed(09.6875,QstateIM(1)) then
				char1IM <= "+09.6875";
			elsif QstateIM(1) = to_sfixed(09.7500,QstateIM(1)) then
				char1IM <= "+09.7500";
			elsif QstateIM(1) = to_sfixed(09.8125,QstateIM(1)) then
				char1IM <= "+09.8125";
			elsif QstateIM(1) = to_sfixed(09.8750,QstateIM(1)) then
				char1IM <= "+09.8750";
			elsif QstateIM(1) = to_sfixed(09.9375,QstateIM(1)) then
				char1IM <= "+09.9375";
			elsif QstateIM(1) = to_sfixed(10.0000,QstateIM(1)) then
				char1IM <= "+10.0000";
			elsif QstateIM(1) = to_sfixed(10.0625,QstateIM(1)) then
				char1IM <= "+10.0625";
			elsif QstateIM(1) = to_sfixed(10.1250,QstateIM(1)) then
				char1IM <= "+10.1250";
			elsif QstateIM(1) = to_sfixed(10.1875,QstateIM(1)) then
				char1IM <= "+10.1875";
			elsif QstateIM(1) = to_sfixed(10.2500,QstateIM(1)) then
				char1IM <= "+10.2500";
			elsif QstateIM(1) = to_sfixed(10.3125,QstateIM(1)) then
				char1IM <= "+10.3125";
			elsif QstateIM(1) = to_sfixed(10.3750,QstateIM(1)) then
				char1IM <= "+10.3750";
			elsif QstateIM(1) = to_sfixed(10.4375,QstateIM(1)) then
				char1IM <= "+10.4375";
			elsif QstateIM(1) = to_sfixed(10.5000,QstateIM(1)) then
				char1IM <= "+10.5000";
			elsif QstateIM(1) = to_sfixed(10.5625,QstateIM(1)) then
				char1IM <= "+10.5625";
			elsif QstateIM(1) = to_sfixed(10.6250,QstateIM(1)) then
				char1IM <= "+10.6250";
			elsif QstateIM(1) = to_sfixed(10.6875,QstateIM(1)) then
				char1IM <= "+10.6875";
			elsif QstateIM(1) = to_sfixed(10.7500,QstateIM(1)) then
				char1IM <= "+10.7500";
			elsif QstateIM(1) = to_sfixed(10.8125,QstateIM(1)) then
				char1IM <= "+10.8125";
			elsif QstateIM(1) = to_sfixed(10.8750,QstateIM(1)) then
				char1IM <= "+10.8750";
			elsif QstateIM(1) = to_sfixed(10.9375,QstateIM(1)) then
				char1IM <= "+10.9375";
			elsif QstateIM(1) = to_sfixed(11.0000,QstateIM(1)) then
				char1IM <= "+11.0000";
			elsif QstateIM(1) = to_sfixed(11.0625,QstateIM(1)) then
				char1IM <= "+11.0625";
			elsif QstateIM(1) = to_sfixed(11.1250,QstateIM(1)) then
				char1IM <= "+11.1250";
			elsif QstateIM(1) = to_sfixed(11.1875,QstateIM(1)) then
				char1IM <= "+11.1875";
			elsif QstateIM(1) = to_sfixed(11.2500,QstateIM(1)) then
				char1IM <= "+11.2500";
			elsif QstateIM(1) = to_sfixed(11.3125,QstateIM(1)) then
				char1IM <= "+11.3125";
			elsif QstateIM(1) = to_sfixed(11.3750,QstateIM(1)) then
				char1IM <= "+11.3750";
			elsif QstateIM(1) = to_sfixed(11.4375,QstateIM(1)) then
				char1IM <= "+11.4375";
			elsif QstateIM(1) = to_sfixed(11.5000,QstateIM(1)) then
				char1IM <= "+11.5000";
			elsif QstateIM(1) = to_sfixed(11.5625,QstateIM(1)) then
				char1IM <= "+11.5625";
			elsif QstateIM(1) = to_sfixed(11.6250,QstateIM(1)) then
				char1IM <= "+11.6250";
			elsif QstateIM(1) = to_sfixed(11.6875,QstateIM(1)) then
				char1IM <= "+11.6875";
			elsif QstateIM(1) = to_sfixed(11.7500,QstateIM(1)) then
				char1IM <= "+11.7500";
			elsif QstateIM(1) = to_sfixed(11.8125,QstateIM(1)) then
				char1IM <= "+11.8125";
			elsif QstateIM(1) = to_sfixed(11.8750,QstateIM(1)) then
				char1IM <= "+11.8750";
			elsif QstateIM(1) = to_sfixed(11.9375,QstateIM(1)) then
				char1IM <= "+11.9375";
			elsif QstateIM(1) = to_sfixed(12.0000,QstateIM(1)) then
				char1IM <= "+12.0000";
			elsif QstateIM(1) = to_sfixed(12.0625,QstateIM(1)) then
				char1IM <= "+12.0625";
			elsif QstateIM(1) = to_sfixed(12.1250,QstateIM(1)) then
				char1IM <= "+12.1250";
			elsif QstateIM(1) = to_sfixed(12.1875,QstateIM(1)) then
				char1IM <= "+12.1875";
			elsif QstateIM(1) = to_sfixed(12.2500,QstateIM(1)) then
				char1IM <= "+12.2500";
			elsif QstateIM(1) = to_sfixed(12.3125,QstateIM(1)) then
				char1IM <= "+12.3125";
			elsif QstateIM(1) = to_sfixed(12.3750,QstateIM(1)) then
				char1IM <= "+12.3750";
			elsif QstateIM(1) = to_sfixed(12.4375,QstateIM(1)) then
				char1IM <= "+12.4375";
			elsif QstateIM(1) = to_sfixed(12.5000,QstateIM(1)) then
				char1IM <= "+12.5000";
			elsif QstateIM(1) = to_sfixed(12.5625,QstateIM(1)) then
				char1IM <= "+12.5625";
			elsif QstateIM(1) = to_sfixed(12.6250,QstateIM(1)) then
				char1IM <= "+12.6250";
			elsif QstateIM(1) = to_sfixed(12.6875,QstateIM(1)) then
				char1IM <= "+12.6875";
			elsif QstateIM(1) = to_sfixed(12.7500,QstateIM(1)) then
				char1IM <= "+12.7500";
			elsif QstateIM(1) = to_sfixed(12.8125,QstateIM(1)) then
				char1IM <= "+12.8125";
			elsif QstateIM(1) = to_sfixed(12.8750,QstateIM(1)) then
				char1IM <= "+12.8750";
			elsif QstateIM(1) = to_sfixed(12.9375,QstateIM(1)) then
				char1IM <= "+12.9375";
			elsif QstateIM(1) = to_sfixed(13.0000,QstateIM(1)) then
				char1IM <= "+13.0000";
			elsif QstateIM(1) = to_sfixed(13.0625,QstateIM(1)) then
				char1IM <= "+13.0625";
			elsif QstateIM(1) = to_sfixed(13.1250,QstateIM(1)) then
				char1IM <= "+13.1250";
			elsif QstateIM(1) = to_sfixed(13.1875,QstateIM(1)) then
				char1IM <= "+13.1875";
			elsif QstateIM(1) = to_sfixed(13.2500,QstateIM(1)) then
				char1IM <= "+13.2500";
			elsif QstateIM(1) = to_sfixed(13.3125,QstateIM(1)) then
				char1IM <= "+13.3125";
			elsif QstateIM(1) = to_sfixed(13.3750,QstateIM(1)) then
				char1IM <= "+13.3750";
			elsif QstateIM(1) = to_sfixed(13.4375,QstateIM(1)) then
				char1IM <= "+13.4375";
			elsif QstateIM(1) = to_sfixed(13.5000,QstateIM(1)) then
				char1IM <= "+13.5000";
			elsif QstateIM(1) = to_sfixed(13.5625,QstateIM(1)) then
				char1IM <= "+13.5625";
			elsif QstateIM(1) = to_sfixed(13.6250,QstateIM(1)) then
				char1IM <= "+13.6250";
			elsif QstateIM(1) = to_sfixed(13.6875,QstateIM(1)) then
				char1IM <= "+13.6875";
			elsif QstateIM(1) = to_sfixed(13.7500,QstateIM(1)) then
				char1IM <= "+13.7500";
			elsif QstateIM(1) = to_sfixed(13.8125,QstateIM(1)) then
				char1IM <= "+13.8125";
			elsif QstateIM(1) = to_sfixed(13.8750,QstateIM(1)) then
				char1IM <= "+13.8750";
			elsif QstateIM(1) = to_sfixed(13.9375,QstateIM(1)) then
				char1IM <= "+13.9375";
			elsif QstateIM(1) = to_sfixed(14.0000,QstateIM(1)) then
				char1IM <= "+14.0000";
			elsif QstateIM(1) = to_sfixed(14.0625,QstateIM(1)) then
				char1IM <= "+14.0625";
			elsif QstateIM(1) = to_sfixed(14.1250,QstateIM(1)) then
				char1IM <= "+14.1250";
			elsif QstateIM(1) = to_sfixed(14.1875,QstateIM(1)) then
				char1IM <= "+14.1875";
			elsif QstateIM(1) = to_sfixed(14.2500,QstateIM(1)) then
				char1IM <= "+14.2500";
			elsif QstateIM(1) = to_sfixed(14.3125,QstateIM(1)) then
				char1IM <= "+14.3125";
			elsif QstateIM(1) = to_sfixed(14.3750,QstateIM(1)) then
				char1IM <= "+14.3750";
			elsif QstateIM(1) = to_sfixed(14.4375,QstateIM(1)) then
				char1IM <= "+14.4375";
			elsif QstateIM(1) = to_sfixed(14.5000,QstateIM(1)) then
				char1IM <= "+14.5000";
			elsif QstateIM(1) = to_sfixed(14.5625,QstateIM(1)) then
				char1IM <= "+14.5625";
			elsif QstateIM(1) = to_sfixed(14.6250,QstateIM(1)) then
				char1IM <= "+14.6250";
			elsif QstateIM(1) = to_sfixed(14.6875,QstateIM(1)) then
				char1IM <= "+14.6875";
			elsif QstateIM(1) = to_sfixed(14.7500,QstateIM(1)) then
				char1IM <= "+14.7500";
			elsif QstateIM(1) = to_sfixed(14.8125,QstateIM(1)) then
				char1IM <= "+14.8125";
			elsif QstateIM(1) = to_sfixed(14.8750,QstateIM(1)) then
				char1IM <= "+14.8750";
			elsif QstateIM(1) = to_sfixed(14.9375,QstateIM(1)) then
				char1IM <= "+14.9375";
			elsif QstateIM(1) = to_sfixed(15.0000,QstateIM(1)) then
				char1IM <= "+15.0000";
			elsif QstateIM(1) = to_sfixed(15.0625,QstateIM(1)) then
				char1IM <= "+15.0625";
			elsif QstateIM(1) = to_sfixed(15.1250,QstateIM(1)) then
				char1IM <= "+15.1250";
			elsif QstateIM(1) = to_sfixed(15.1875,QstateIM(1)) then
				char1IM <= "+15.1875";
			elsif QstateIM(1) = to_sfixed(15.2500,QstateIM(1)) then
				char1IM <= "+15.2500";
			elsif QstateIM(1) = to_sfixed(15.3125,QstateIM(1)) then
				char1IM <= "+15.3125";
			elsif QstateIM(1) = to_sfixed(15.3750,QstateIM(1)) then
				char1IM <= "+15.3750";
			elsif QstateIM(1) = to_sfixed(15.4375,QstateIM(1)) then
				char1IM <= "+15.4375";
			elsif QstateIM(1) = to_sfixed(15.5000,QstateIM(1)) then
				char1IM <= "+15.5000";
			elsif QstateIM(1) = to_sfixed(15.5625,QstateIM(1)) then
				char1IM <= "+15.5625";
			elsif QstateIM(1) = to_sfixed(15.6250,QstateIM(1)) then
				char1IM <= "+15.6250";
			elsif QstateIM(1) = to_sfixed(15.6875,QstateIM(1)) then
				char1IM <= "+15.6875";
			elsif QstateIM(1) = to_sfixed(15.7500,QstateIM(1)) then
				char1IM <= "+15.7500";
			elsif QstateIM(1) = to_sfixed(15.8125,QstateIM(1)) then
				char1IM <= "+15.8125";
			elsif QstateIM(1) = to_sfixed(15.8750,QstateIM(1)) then
				char1IM <= "+15.8750";
			elsif QstateIM(1) = to_sfixed(15.9375,QstateIM(1)) then
				char1IM <= "+15.9375";
			end if;
			if QstateRE(2) = to_sfixed(-15.9375,QstateRE(2)) then
				char2RE <= "-15.9375";
			elsif QstateRE(2) = to_sfixed(-15.8750,QstateRE(2)) then
				char2RE <= "-15.8750";
			elsif QstateRE(2) = to_sfixed(-15.8125,QstateRE(2)) then
				char2RE <= "-15.8125";
			elsif QstateRE(2) = to_sfixed(-15.7500,QstateRE(2)) then
				char2RE <= "-15.7500";
			elsif QstateRE(2) = to_sfixed(-15.6875,QstateRE(2)) then
				char2RE <= "-15.6875";
			elsif QstateRE(2) = to_sfixed(-15.6250,QstateRE(2)) then
				char2RE <= "-15.6250";
			elsif QstateRE(2) = to_sfixed(-15.5625,QstateRE(2)) then
				char2RE <= "-15.5625";
			elsif QstateRE(2) = to_sfixed(-15.5000,QstateRE(2)) then
				char2RE <= "-15.5000";
			elsif QstateRE(2) = to_sfixed(-15.4375,QstateRE(2)) then
				char2RE <= "-15.4375";
			elsif QstateRE(2) = to_sfixed(-15.3750,QstateRE(2)) then
				char2RE <= "-15.3750";
			elsif QstateRE(2) = to_sfixed(-15.3125,QstateRE(2)) then
				char2RE <= "-15.3125";
			elsif QstateRE(2) = to_sfixed(-15.2500,QstateRE(2)) then
				char2RE <= "-15.2500";
			elsif QstateRE(2) = to_sfixed(-15.1875,QstateRE(2)) then
				char2RE <= "-15.1875";
			elsif QstateRE(2) = to_sfixed(-15.1250,QstateRE(2)) then
				char2RE <= "-15.1250";
			elsif QstateRE(2) = to_sfixed(-15.0625,QstateRE(2)) then
				char2RE <= "-15.0625";
			elsif QstateRE(2) = to_sfixed(-15.0000,QstateRE(2)) then
				char2RE <= "-15.0000";
			elsif QstateRE(2) = to_sfixed(-14.9375,QstateRE(2)) then
				char2RE <= "-14.9375";
			elsif QstateRE(2) = to_sfixed(-14.8750,QstateRE(2)) then
				char2RE <= "-14.8750";
			elsif QstateRE(2) = to_sfixed(-14.8125,QstateRE(2)) then
				char2RE <= "-14.8125";
			elsif QstateRE(2) = to_sfixed(-14.7500,QstateRE(2)) then
				char2RE <= "-14.7500";
			elsif QstateRE(2) = to_sfixed(-14.6875,QstateRE(2)) then
				char2RE <= "-14.6875";
			elsif QstateRE(2) = to_sfixed(-14.6250,QstateRE(2)) then
				char2RE <= "-14.6250";
			elsif QstateRE(2) = to_sfixed(-14.5625,QstateRE(2)) then
				char2RE <= "-14.5625";
			elsif QstateRE(2) = to_sfixed(-14.5000,QstateRE(2)) then
				char2RE <= "-14.5000";
			elsif QstateRE(2) = to_sfixed(-14.4375,QstateRE(2)) then
				char2RE <= "-14.4375";
			elsif QstateRE(2) = to_sfixed(-14.3750,QstateRE(2)) then
				char2RE <= "-14.3750";
			elsif QstateRE(2) = to_sfixed(-14.3125,QstateRE(2)) then
				char2RE <= "-14.3125";
			elsif QstateRE(2) = to_sfixed(-14.2500,QstateRE(2)) then
				char2RE <= "-14.2500";
			elsif QstateRE(2) = to_sfixed(-14.1875,QstateRE(2)) then
				char2RE <= "-14.1875";
			elsif QstateRE(2) = to_sfixed(-14.1250,QstateRE(2)) then
				char2RE <= "-14.1250";
			elsif QstateRE(2) = to_sfixed(-14.0625,QstateRE(2)) then
				char2RE <= "-14.0625";
			elsif QstateRE(2) = to_sfixed(-14.0000,QstateRE(2)) then
				char2RE <= "-14.0000";
			elsif QstateRE(2) = to_sfixed(-13.9375,QstateRE(2)) then
				char2RE <= "-13.9375";
			elsif QstateRE(2) = to_sfixed(-13.8750,QstateRE(2)) then
				char2RE <= "-13.8750";
			elsif QstateRE(2) = to_sfixed(-13.8125,QstateRE(2)) then
				char2RE <= "-13.8125";
			elsif QstateRE(2) = to_sfixed(-13.7500,QstateRE(2)) then
				char2RE <= "-13.7500";
			elsif QstateRE(2) = to_sfixed(-13.6875,QstateRE(2)) then
				char2RE <= "-13.6875";
			elsif QstateRE(2) = to_sfixed(-13.6250,QstateRE(2)) then
				char2RE <= "-13.6250";
			elsif QstateRE(2) = to_sfixed(-13.5625,QstateRE(2)) then
				char2RE <= "-13.5625";
			elsif QstateRE(2) = to_sfixed(-13.5000,QstateRE(2)) then
				char2RE <= "-13.5000";
			elsif QstateRE(2) = to_sfixed(-13.4375,QstateRE(2)) then
				char2RE <= "-13.4375";
			elsif QstateRE(2) = to_sfixed(-13.3750,QstateRE(2)) then
				char2RE <= "-13.3750";
			elsif QstateRE(2) = to_sfixed(-13.3125,QstateRE(2)) then
				char2RE <= "-13.3125";
			elsif QstateRE(2) = to_sfixed(-13.2500,QstateRE(2)) then
				char2RE <= "-13.2500";
			elsif QstateRE(2) = to_sfixed(-13.1875,QstateRE(2)) then
				char2RE <= "-13.1875";
			elsif QstateRE(2) = to_sfixed(-13.1250,QstateRE(2)) then
				char2RE <= "-13.1250";
			elsif QstateRE(2) = to_sfixed(-13.0625,QstateRE(2)) then
				char2RE <= "-13.0625";
			elsif QstateRE(2) = to_sfixed(-13.0000,QstateRE(2)) then
				char2RE <= "-13.0000";
			elsif QstateRE(2) = to_sfixed(-12.9375,QstateRE(2)) then
				char2RE <= "-12.9375";
			elsif QstateRE(2) = to_sfixed(-12.8750,QstateRE(2)) then
				char2RE <= "-12.8750";
			elsif QstateRE(2) = to_sfixed(-12.8125,QstateRE(2)) then
				char2RE <= "-12.8125";
			elsif QstateRE(2) = to_sfixed(-12.7500,QstateRE(2)) then
				char2RE <= "-12.7500";
			elsif QstateRE(2) = to_sfixed(-12.6875,QstateRE(2)) then
				char2RE <= "-12.6875";
			elsif QstateRE(2) = to_sfixed(-12.6250,QstateRE(2)) then
				char2RE <= "-12.6250";
			elsif QstateRE(2) = to_sfixed(-12.5625,QstateRE(2)) then
				char2RE <= "-12.5625";
			elsif QstateRE(2) = to_sfixed(-12.5000,QstateRE(2)) then
				char2RE <= "-12.5000";
			elsif QstateRE(2) = to_sfixed(-12.4375,QstateRE(2)) then
				char2RE <= "-12.4375";
			elsif QstateRE(2) = to_sfixed(-12.3750,QstateRE(2)) then
				char2RE <= "-12.3750";
			elsif QstateRE(2) = to_sfixed(-12.3125,QstateRE(2)) then
				char2RE <= "-12.3125";
			elsif QstateRE(2) = to_sfixed(-12.2500,QstateRE(2)) then
				char2RE <= "-12.2500";
			elsif QstateRE(2) = to_sfixed(-12.1875,QstateRE(2)) then
				char2RE <= "-12.1875";
			elsif QstateRE(2) = to_sfixed(-12.1250,QstateRE(2)) then
				char2RE <= "-12.1250";
			elsif QstateRE(2) = to_sfixed(-12.0625,QstateRE(2)) then
				char2RE <= "-12.0625";
			elsif QstateRE(2) = to_sfixed(-12.0000,QstateRE(2)) then
				char2RE <= "-12.0000";
			elsif QstateRE(2) = to_sfixed(-11.9375,QstateRE(2)) then
				char2RE <= "-11.9375";
			elsif QstateRE(2) = to_sfixed(-11.8750,QstateRE(2)) then
				char2RE <= "-11.8750";
			elsif QstateRE(2) = to_sfixed(-11.8125,QstateRE(2)) then
				char2RE <= "-11.8125";
			elsif QstateRE(2) = to_sfixed(-11.7500,QstateRE(2)) then
				char2RE <= "-11.7500";
			elsif QstateRE(2) = to_sfixed(-11.6875,QstateRE(2)) then
				char2RE <= "-11.6875";
			elsif QstateRE(2) = to_sfixed(-11.6250,QstateRE(2)) then
				char2RE <= "-11.6250";
			elsif QstateRE(2) = to_sfixed(-11.5625,QstateRE(2)) then
				char2RE <= "-11.5625";
			elsif QstateRE(2) = to_sfixed(-11.5000,QstateRE(2)) then
				char2RE <= "-11.5000";
			elsif QstateRE(2) = to_sfixed(-11.4375,QstateRE(2)) then
				char2RE <= "-11.4375";
			elsif QstateRE(2) = to_sfixed(-11.3750,QstateRE(2)) then
				char2RE <= "-11.3750";
			elsif QstateRE(2) = to_sfixed(-11.3125,QstateRE(2)) then
				char2RE <= "-11.3125";
			elsif QstateRE(2) = to_sfixed(-11.2500,QstateRE(2)) then
				char2RE <= "-11.2500";
			elsif QstateRE(2) = to_sfixed(-11.1875,QstateRE(2)) then
				char2RE <= "-11.1875";
			elsif QstateRE(2) = to_sfixed(-11.1250,QstateRE(2)) then
				char2RE <= "-11.1250";
			elsif QstateRE(2) = to_sfixed(-11.0625,QstateRE(2)) then
				char2RE <= "-11.0625";
			elsif QstateRE(2) = to_sfixed(-11.0000,QstateRE(2)) then
				char2RE <= "-11.0000";
			elsif QstateRE(2) = to_sfixed(-10.9375,QstateRE(2)) then
				char2RE <= "-10.9375";
			elsif QstateRE(2) = to_sfixed(-10.8750,QstateRE(2)) then
				char2RE <= "-10.8750";
			elsif QstateRE(2) = to_sfixed(-10.8125,QstateRE(2)) then
				char2RE <= "-10.8125";
			elsif QstateRE(2) = to_sfixed(-10.7500,QstateRE(2)) then
				char2RE <= "-10.7500";
			elsif QstateRE(2) = to_sfixed(-10.6875,QstateRE(2)) then
				char2RE <= "-10.6875";
			elsif QstateRE(2) = to_sfixed(-10.6250,QstateRE(2)) then
				char2RE <= "-10.6250";
			elsif QstateRE(2) = to_sfixed(-10.5625,QstateRE(2)) then
				char2RE <= "-10.5625";
			elsif QstateRE(2) = to_sfixed(-10.5000,QstateRE(2)) then
				char2RE <= "-10.5000";
			elsif QstateRE(2) = to_sfixed(-10.4375,QstateRE(2)) then
				char2RE <= "-10.4375";
			elsif QstateRE(2) = to_sfixed(-10.3750,QstateRE(2)) then
				char2RE <= "-10.3750";
			elsif QstateRE(2) = to_sfixed(-10.3125,QstateRE(2)) then
				char2RE <= "-10.3125";
			elsif QstateRE(2) = to_sfixed(-10.2500,QstateRE(2)) then
				char2RE <= "-10.2500";
			elsif QstateRE(2) = to_sfixed(-10.1875,QstateRE(2)) then
				char2RE <= "-10.1875";
			elsif QstateRE(2) = to_sfixed(-10.1250,QstateRE(2)) then
				char2RE <= "-10.1250";
			elsif QstateRE(2) = to_sfixed(-10.0625,QstateRE(2)) then
				char2RE <= "-10.0625";
			elsif QstateRE(2) = to_sfixed(-10.0000,QstateRE(2)) then
				char2RE <= "-10.0000";
			elsif QstateRE(2) = to_sfixed(-9.9375,QstateRE(2)) then
				char2RE <= "--9.9375";
			elsif QstateRE(2) = to_sfixed(-9.8750,QstateRE(2)) then
				char2RE <= "--9.8750";
			elsif QstateRE(2) = to_sfixed(-9.8125,QstateRE(2)) then
				char2RE <= "--9.8125";
			elsif QstateRE(2) = to_sfixed(-9.7500,QstateRE(2)) then
				char2RE <= "--9.7500";
			elsif QstateRE(2) = to_sfixed(-9.6875,QstateRE(2)) then
				char2RE <= "--9.6875";
			elsif QstateRE(2) = to_sfixed(-9.6250,QstateRE(2)) then
				char2RE <= "--9.6250";
			elsif QstateRE(2) = to_sfixed(-9.5625,QstateRE(2)) then
				char2RE <= "--9.5625";
			elsif QstateRE(2) = to_sfixed(-9.5000,QstateRE(2)) then
				char2RE <= "--9.5000";
			elsif QstateRE(2) = to_sfixed(-9.4375,QstateRE(2)) then
				char2RE <= "--9.4375";
			elsif QstateRE(2) = to_sfixed(-9.3750,QstateRE(2)) then
				char2RE <= "--9.3750";
			elsif QstateRE(2) = to_sfixed(-9.3125,QstateRE(2)) then
				char2RE <= "--9.3125";
			elsif QstateRE(2) = to_sfixed(-9.2500,QstateRE(2)) then
				char2RE <= "--9.2500";
			elsif QstateRE(2) = to_sfixed(-9.1875,QstateRE(2)) then
				char2RE <= "--9.1875";
			elsif QstateRE(2) = to_sfixed(-9.1250,QstateRE(2)) then
				char2RE <= "--9.1250";
			elsif QstateRE(2) = to_sfixed(-9.0625,QstateRE(2)) then
				char2RE <= "--9.0625";
			elsif QstateRE(2) = to_sfixed(-9.0000,QstateRE(2)) then
				char2RE <= "--9.0000";
			elsif QstateRE(2) = to_sfixed(-8.9375,QstateRE(2)) then
				char2RE <= "--8.9375";
			elsif QstateRE(2) = to_sfixed(-8.8750,QstateRE(2)) then
				char2RE <= "--8.8750";
			elsif QstateRE(2) = to_sfixed(-8.8125,QstateRE(2)) then
				char2RE <= "--8.8125";
			elsif QstateRE(2) = to_sfixed(-8.7500,QstateRE(2)) then
				char2RE <= "--8.7500";
			elsif QstateRE(2) = to_sfixed(-8.6875,QstateRE(2)) then
				char2RE <= "--8.6875";
			elsif QstateRE(2) = to_sfixed(-8.6250,QstateRE(2)) then
				char2RE <= "--8.6250";
			elsif QstateRE(2) = to_sfixed(-8.5625,QstateRE(2)) then
				char2RE <= "--8.5625";
			elsif QstateRE(2) = to_sfixed(-8.5000,QstateRE(2)) then
				char2RE <= "--8.5000";
			elsif QstateRE(2) = to_sfixed(-8.4375,QstateRE(2)) then
				char2RE <= "--8.4375";
			elsif QstateRE(2) = to_sfixed(-8.3750,QstateRE(2)) then
				char2RE <= "--8.3750";
			elsif QstateRE(2) = to_sfixed(-8.3125,QstateRE(2)) then
				char2RE <= "--8.3125";
			elsif QstateRE(2) = to_sfixed(-8.2500,QstateRE(2)) then
				char2RE <= "--8.2500";
			elsif QstateRE(2) = to_sfixed(-8.1875,QstateRE(2)) then
				char2RE <= "--8.1875";
			elsif QstateRE(2) = to_sfixed(-8.1250,QstateRE(2)) then
				char2RE <= "--8.1250";
			elsif QstateRE(2) = to_sfixed(-8.0625,QstateRE(2)) then
				char2RE <= "--8.0625";
			elsif QstateRE(2) = to_sfixed(-8.0000,QstateRE(2)) then
				char2RE <= "--8.0000";
			elsif QstateRE(2) = to_sfixed(-7.9375,QstateRE(2)) then
				char2RE <= "--7.9375";
			elsif QstateRE(2) = to_sfixed(-7.8750,QstateRE(2)) then
				char2RE <= "--7.8750";
			elsif QstateRE(2) = to_sfixed(-7.8125,QstateRE(2)) then
				char2RE <= "--7.8125";
			elsif QstateRE(2) = to_sfixed(-7.7500,QstateRE(2)) then
				char2RE <= "--7.7500";
			elsif QstateRE(2) = to_sfixed(-7.6875,QstateRE(2)) then
				char2RE <= "--7.6875";
			elsif QstateRE(2) = to_sfixed(-7.6250,QstateRE(2)) then
				char2RE <= "--7.6250";
			elsif QstateRE(2) = to_sfixed(-7.5625,QstateRE(2)) then
				char2RE <= "--7.5625";
			elsif QstateRE(2) = to_sfixed(-7.5000,QstateRE(2)) then
				char2RE <= "--7.5000";
			elsif QstateRE(2) = to_sfixed(-7.4375,QstateRE(2)) then
				char2RE <= "--7.4375";
			elsif QstateRE(2) = to_sfixed(-7.3750,QstateRE(2)) then
				char2RE <= "--7.3750";
			elsif QstateRE(2) = to_sfixed(-7.3125,QstateRE(2)) then
				char2RE <= "--7.3125";
			elsif QstateRE(2) = to_sfixed(-7.2500,QstateRE(2)) then
				char2RE <= "--7.2500";
			elsif QstateRE(2) = to_sfixed(-7.1875,QstateRE(2)) then
				char2RE <= "--7.1875";
			elsif QstateRE(2) = to_sfixed(-7.1250,QstateRE(2)) then
				char2RE <= "--7.1250";
			elsif QstateRE(2) = to_sfixed(-7.0625,QstateRE(2)) then
				char2RE <= "--7.0625";
			elsif QstateRE(2) = to_sfixed(-7.0000,QstateRE(2)) then
				char2RE <= "--7.0000";
			elsif QstateRE(2) = to_sfixed(-6.9375,QstateRE(2)) then
				char2RE <= "--6.9375";
			elsif QstateRE(2) = to_sfixed(-6.8750,QstateRE(2)) then
				char2RE <= "--6.8750";
			elsif QstateRE(2) = to_sfixed(-6.8125,QstateRE(2)) then
				char2RE <= "--6.8125";
			elsif QstateRE(2) = to_sfixed(-6.7500,QstateRE(2)) then
				char2RE <= "--6.7500";
			elsif QstateRE(2) = to_sfixed(-6.6875,QstateRE(2)) then
				char2RE <= "--6.6875";
			elsif QstateRE(2) = to_sfixed(-6.6250,QstateRE(2)) then
				char2RE <= "--6.6250";
			elsif QstateRE(2) = to_sfixed(-6.5625,QstateRE(2)) then
				char2RE <= "--6.5625";
			elsif QstateRE(2) = to_sfixed(-6.5000,QstateRE(2)) then
				char2RE <= "--6.5000";
			elsif QstateRE(2) = to_sfixed(-6.4375,QstateRE(2)) then
				char2RE <= "--6.4375";
			elsif QstateRE(2) = to_sfixed(-6.3750,QstateRE(2)) then
				char2RE <= "--6.3750";
			elsif QstateRE(2) = to_sfixed(-6.3125,QstateRE(2)) then
				char2RE <= "--6.3125";
			elsif QstateRE(2) = to_sfixed(-6.2500,QstateRE(2)) then
				char2RE <= "--6.2500";
			elsif QstateRE(2) = to_sfixed(-6.1875,QstateRE(2)) then
				char2RE <= "--6.1875";
			elsif QstateRE(2) = to_sfixed(-6.1250,QstateRE(2)) then
				char2RE <= "--6.1250";
			elsif QstateRE(2) = to_sfixed(-6.0625,QstateRE(2)) then
				char2RE <= "--6.0625";
			elsif QstateRE(2) = to_sfixed(-6.0000,QstateRE(2)) then
				char2RE <= "--6.0000";
			elsif QstateRE(2) = to_sfixed(-5.9375,QstateRE(2)) then
				char2RE <= "--5.9375";
			elsif QstateRE(2) = to_sfixed(-5.8750,QstateRE(2)) then
				char2RE <= "--5.8750";
			elsif QstateRE(2) = to_sfixed(-5.8125,QstateRE(2)) then
				char2RE <= "--5.8125";
			elsif QstateRE(2) = to_sfixed(-5.7500,QstateRE(2)) then
				char2RE <= "--5.7500";
			elsif QstateRE(2) = to_sfixed(-5.6875,QstateRE(2)) then
				char2RE <= "--5.6875";
			elsif QstateRE(2) = to_sfixed(-5.6250,QstateRE(2)) then
				char2RE <= "--5.6250";
			elsif QstateRE(2) = to_sfixed(-5.5625,QstateRE(2)) then
				char2RE <= "--5.5625";
			elsif QstateRE(2) = to_sfixed(-5.5000,QstateRE(2)) then
				char2RE <= "--5.5000";
			elsif QstateRE(2) = to_sfixed(-5.4375,QstateRE(2)) then
				char2RE <= "--5.4375";
			elsif QstateRE(2) = to_sfixed(-5.3750,QstateRE(2)) then
				char2RE <= "--5.3750";
			elsif QstateRE(2) = to_sfixed(-5.3125,QstateRE(2)) then
				char2RE <= "--5.3125";
			elsif QstateRE(2) = to_sfixed(-5.2500,QstateRE(2)) then
				char2RE <= "--5.2500";
			elsif QstateRE(2) = to_sfixed(-5.1875,QstateRE(2)) then
				char2RE <= "--5.1875";
			elsif QstateRE(2) = to_sfixed(-5.1250,QstateRE(2)) then
				char2RE <= "--5.1250";
			elsif QstateRE(2) = to_sfixed(-5.0625,QstateRE(2)) then
				char2RE <= "--5.0625";
			elsif QstateRE(2) = to_sfixed(-5.0000,QstateRE(2)) then
				char2RE <= "--5.0000";
			elsif QstateRE(2) = to_sfixed(-4.9375,QstateRE(2)) then
				char2RE <= "--4.9375";
			elsif QstateRE(2) = to_sfixed(-4.8750,QstateRE(2)) then
				char2RE <= "--4.8750";
			elsif QstateRE(2) = to_sfixed(-4.8125,QstateRE(2)) then
				char2RE <= "--4.8125";
			elsif QstateRE(2) = to_sfixed(-4.7500,QstateRE(2)) then
				char2RE <= "--4.7500";
			elsif QstateRE(2) = to_sfixed(-4.6875,QstateRE(2)) then
				char2RE <= "--4.6875";
			elsif QstateRE(2) = to_sfixed(-4.6250,QstateRE(2)) then
				char2RE <= "--4.6250";
			elsif QstateRE(2) = to_sfixed(-4.5625,QstateRE(2)) then
				char2RE <= "--4.5625";
			elsif QstateRE(2) = to_sfixed(-4.5000,QstateRE(2)) then
				char2RE <= "--4.5000";
			elsif QstateRE(2) = to_sfixed(-4.4375,QstateRE(2)) then
				char2RE <= "--4.4375";
			elsif QstateRE(2) = to_sfixed(-4.3750,QstateRE(2)) then
				char2RE <= "--4.3750";
			elsif QstateRE(2) = to_sfixed(-4.3125,QstateRE(2)) then
				char2RE <= "--4.3125";
			elsif QstateRE(2) = to_sfixed(-4.2500,QstateRE(2)) then
				char2RE <= "--4.2500";
			elsif QstateRE(2) = to_sfixed(-4.1875,QstateRE(2)) then
				char2RE <= "--4.1875";
			elsif QstateRE(2) = to_sfixed(-4.1250,QstateRE(2)) then
				char2RE <= "--4.1250";
			elsif QstateRE(2) = to_sfixed(-4.0625,QstateRE(2)) then
				char2RE <= "--4.0625";
			elsif QstateRE(2) = to_sfixed(-4.0000,QstateRE(2)) then
				char2RE <= "--4.0000";
			elsif QstateRE(2) = to_sfixed(-3.9375,QstateRE(2)) then
				char2RE <= "--3.9375";
			elsif QstateRE(2) = to_sfixed(-3.8750,QstateRE(2)) then
				char2RE <= "--3.8750";
			elsif QstateRE(2) = to_sfixed(-3.8125,QstateRE(2)) then
				char2RE <= "--3.8125";
			elsif QstateRE(2) = to_sfixed(-3.7500,QstateRE(2)) then
				char2RE <= "--3.7500";
			elsif QstateRE(2) = to_sfixed(-3.6875,QstateRE(2)) then
				char2RE <= "--3.6875";
			elsif QstateRE(2) = to_sfixed(-3.6250,QstateRE(2)) then
				char2RE <= "--3.6250";
			elsif QstateRE(2) = to_sfixed(-3.5625,QstateRE(2)) then
				char2RE <= "--3.5625";
			elsif QstateRE(2) = to_sfixed(-3.5000,QstateRE(2)) then
				char2RE <= "--3.5000";
			elsif QstateRE(2) = to_sfixed(-3.4375,QstateRE(2)) then
				char2RE <= "--3.4375";
			elsif QstateRE(2) = to_sfixed(-3.3750,QstateRE(2)) then
				char2RE <= "--3.3750";
			elsif QstateRE(2) = to_sfixed(-3.3125,QstateRE(2)) then
				char2RE <= "--3.3125";
			elsif QstateRE(2) = to_sfixed(-3.2500,QstateRE(2)) then
				char2RE <= "--3.2500";
			elsif QstateRE(2) = to_sfixed(-3.1875,QstateRE(2)) then
				char2RE <= "--3.1875";
			elsif QstateRE(2) = to_sfixed(-3.1250,QstateRE(2)) then
				char2RE <= "--3.1250";
			elsif QstateRE(2) = to_sfixed(-3.0625,QstateRE(2)) then
				char2RE <= "--3.0625";
			elsif QstateRE(2) = to_sfixed(-3.0000,QstateRE(2)) then
				char2RE <= "--3.0000";
			elsif QstateRE(2) = to_sfixed(-2.9375,QstateRE(2)) then
				char2RE <= "--2.9375";
			elsif QstateRE(2) = to_sfixed(-2.8750,QstateRE(2)) then
				char2RE <= "--2.8750";
			elsif QstateRE(2) = to_sfixed(-2.8125,QstateRE(2)) then
				char2RE <= "--2.8125";
			elsif QstateRE(2) = to_sfixed(-2.7500,QstateRE(2)) then
				char2RE <= "--2.7500";
			elsif QstateRE(2) = to_sfixed(-2.6875,QstateRE(2)) then
				char2RE <= "--2.6875";
			elsif QstateRE(2) = to_sfixed(-2.6250,QstateRE(2)) then
				char2RE <= "--2.6250";
			elsif QstateRE(2) = to_sfixed(-2.5625,QstateRE(2)) then
				char2RE <= "--2.5625";
			elsif QstateRE(2) = to_sfixed(-2.5000,QstateRE(2)) then
				char2RE <= "--2.5000";
			elsif QstateRE(2) = to_sfixed(-2.4375,QstateRE(2)) then
				char2RE <= "--2.4375";
			elsif QstateRE(2) = to_sfixed(-2.3750,QstateRE(2)) then
				char2RE <= "--2.3750";
			elsif QstateRE(2) = to_sfixed(-2.3125,QstateRE(2)) then
				char2RE <= "--2.3125";
			elsif QstateRE(2) = to_sfixed(-2.2500,QstateRE(2)) then
				char2RE <= "--2.2500";
			elsif QstateRE(2) = to_sfixed(-2.1875,QstateRE(2)) then
				char2RE <= "--2.1875";
			elsif QstateRE(2) = to_sfixed(-2.1250,QstateRE(2)) then
				char2RE <= "--2.1250";
			elsif QstateRE(2) = to_sfixed(-2.0625,QstateRE(2)) then
				char2RE <= "--2.0625";
			elsif QstateRE(2) = to_sfixed(-2.0000,QstateRE(2)) then
				char2RE <= "--2.0000";
			elsif QstateRE(2) = to_sfixed(-1.9375,QstateRE(2)) then
				char2RE <= "--1.9375";
			elsif QstateRE(2) = to_sfixed(-1.8750,QstateRE(2)) then
				char2RE <= "--1.8750";
			elsif QstateRE(2) = to_sfixed(-1.8125,QstateRE(2)) then
				char2RE <= "--1.8125";
			elsif QstateRE(2) = to_sfixed(-1.7500,QstateRE(2)) then
				char2RE <= "--1.7500";
			elsif QstateRE(2) = to_sfixed(-1.6875,QstateRE(2)) then
				char2RE <= "--1.6875";
			elsif QstateRE(2) = to_sfixed(-1.6250,QstateRE(2)) then
				char2RE <= "--1.6250";
			elsif QstateRE(2) = to_sfixed(-1.5625,QstateRE(2)) then
				char2RE <= "--1.5625";
			elsif QstateRE(2) = to_sfixed(-1.5000,QstateRE(2)) then
				char2RE <= "--1.5000";
			elsif QstateRE(2) = to_sfixed(-1.4375,QstateRE(2)) then
				char2RE <= "--1.4375";
			elsif QstateRE(2) = to_sfixed(-1.3750,QstateRE(2)) then
				char2RE <= "--1.3750";
			elsif QstateRE(2) = to_sfixed(-1.3125,QstateRE(2)) then
				char2RE <= "--1.3125";
			elsif QstateRE(2) = to_sfixed(-1.2500,QstateRE(2)) then
				char2RE <= "--1.2500";
			elsif QstateRE(2) = to_sfixed(-1.1875,QstateRE(2)) then
				char2RE <= "--1.1875";
			elsif QstateRE(2) = to_sfixed(-1.1250,QstateRE(2)) then
				char2RE <= "--1.1250";
			elsif QstateRE(2) = to_sfixed(-1.0625,QstateRE(2)) then
				char2RE <= "--1.0625";
			elsif QstateRE(2) = to_sfixed(-1.0000,QstateRE(2)) then
				char2RE <= "--1.0000";
			elsif QstateRE(2) = to_sfixed(-0.9375,QstateRE(2)) then
				char2RE <= "--0.9375";
			elsif QstateRE(2) = to_sfixed(-0.8750,QstateRE(2)) then
				char2RE <= "--0.8750";
			elsif QstateRE(2) = to_sfixed(-0.8125,QstateRE(2)) then
				char2RE <= "--0.8125";
			elsif QstateRE(2) = to_sfixed(-0.7500,QstateRE(2)) then
				char2RE <= "--0.7500";
			elsif QstateRE(2) = to_sfixed(-0.6875,QstateRE(2)) then
				char2RE <= "--0.6875";
			elsif QstateRE(2) = to_sfixed(-0.6250,QstateRE(2)) then
				char2RE <= "--0.6250";
			elsif QstateRE(2) = to_sfixed(-0.5625,QstateRE(2)) then
				char2RE <= "--0.5625";
			elsif QstateRE(2) = to_sfixed(-0.5000,QstateRE(2)) then
				char2RE <= "--0.5000";
			elsif QstateRE(2) = to_sfixed(-0.4375,QstateRE(2)) then
				char2RE <= "--0.4375";
			elsif QstateRE(2) = to_sfixed(-0.3750,QstateRE(2)) then
				char2RE <= "--0.3750";
			elsif QstateRE(2) = to_sfixed(-0.3125,QstateRE(2)) then
				char2RE <= "--0.3125";
			elsif QstateRE(2) = to_sfixed(-0.2500,QstateRE(2)) then
				char2RE <= "--0.2500";
			elsif QstateRE(2) = to_sfixed(-0.1875,QstateRE(2)) then
				char2RE <= "--0.1875";
			elsif QstateRE(2) = to_sfixed(-0.1250,QstateRE(2)) then
				char2RE <= "--0.1250";
			elsif QstateRE(2) = to_sfixed(-0.0625,QstateRE(2)) then
				char2RE <= "--0.0625";
			elsif QstateRE(2) = to_sfixed(00.0000,QstateRE(2)) then
				char2RE <= "+00.0000";
			elsif QstateRE(2) = to_sfixed(00.0625,QstateRE(2)) then
				char2RE <= "+00.0625";
			elsif QstateRE(2) = to_sfixed(00.1250,QstateRE(2)) then
				char2RE <= "+00.1250";
			elsif QstateRE(2) = to_sfixed(00.1875,QstateRE(2)) then
				char2RE <= "+00.1875";
			elsif QstateRE(2) = to_sfixed(00.2500,QstateRE(2)) then
				char2RE <= "+00.2500";
			elsif QstateRE(2) = to_sfixed(00.3125,QstateRE(2)) then
				char2RE <= "+00.3125";
			elsif QstateRE(2) = to_sfixed(00.3750,QstateRE(2)) then
				char2RE <= "+00.3750";
			elsif QstateRE(2) = to_sfixed(00.4375,QstateRE(2)) then
				char2RE <= "+00.4375";
			elsif QstateRE(2) = to_sfixed(00.5000,QstateRE(2)) then
				char2RE <= "+00.5000";
			elsif QstateRE(2) = to_sfixed(00.5625,QstateRE(2)) then
				char2RE <= "+00.5625";
			elsif QstateRE(2) = to_sfixed(00.6250,QstateRE(2)) then
				char2RE <= "+00.6250";
			elsif QstateRE(2) = to_sfixed(00.6875,QstateRE(2)) then
				char2RE <= "+00.6875";
			elsif QstateRE(2) = to_sfixed(00.7500,QstateRE(2)) then
				char2RE <= "+00.7500";
			elsif QstateRE(2) = to_sfixed(00.8125,QstateRE(2)) then
				char2RE <= "+00.8125";
			elsif QstateRE(2) = to_sfixed(00.8750,QstateRE(2)) then
				char2RE <= "+00.8750";
			elsif QstateRE(2) = to_sfixed(00.9375,QstateRE(2)) then
				char2RE <= "+00.9375";
			elsif QstateRE(2) = to_sfixed(01.0000,QstateRE(2)) then
				char2RE <= "+01.0000";
			elsif QstateRE(2) = to_sfixed(01.0625,QstateRE(2)) then
				char2RE <= "+01.0625";
			elsif QstateRE(2) = to_sfixed(01.1250,QstateRE(2)) then
				char2RE <= "+01.1250";
			elsif QstateRE(2) = to_sfixed(01.1875,QstateRE(2)) then
				char2RE <= "+01.1875";
			elsif QstateRE(2) = to_sfixed(01.2500,QstateRE(2)) then
				char2RE <= "+01.2500";
			elsif QstateRE(2) = to_sfixed(01.3125,QstateRE(2)) then
				char2RE <= "+01.3125";
			elsif QstateRE(2) = to_sfixed(01.3750,QstateRE(2)) then
				char2RE <= "+01.3750";
			elsif QstateRE(2) = to_sfixed(01.4375,QstateRE(2)) then
				char2RE <= "+01.4375";
			elsif QstateRE(2) = to_sfixed(01.5000,QstateRE(2)) then
				char2RE <= "+01.5000";
			elsif QstateRE(2) = to_sfixed(01.5625,QstateRE(2)) then
				char2RE <= "+01.5625";
			elsif QstateRE(2) = to_sfixed(01.6250,QstateRE(2)) then
				char2RE <= "+01.6250";
			elsif QstateRE(2) = to_sfixed(01.6875,QstateRE(2)) then
				char2RE <= "+01.6875";
			elsif QstateRE(2) = to_sfixed(01.7500,QstateRE(2)) then
				char2RE <= "+01.7500";
			elsif QstateRE(2) = to_sfixed(01.8125,QstateRE(2)) then
				char2RE <= "+01.8125";
			elsif QstateRE(2) = to_sfixed(01.8750,QstateRE(2)) then
				char2RE <= "+01.8750";
			elsif QstateRE(2) = to_sfixed(01.9375,QstateRE(2)) then
				char2RE <= "+01.9375";
			elsif QstateRE(2) = to_sfixed(02.0000,QstateRE(2)) then
				char2RE <= "+02.0000";
			elsif QstateRE(2) = to_sfixed(02.0625,QstateRE(2)) then
				char2RE <= "+02.0625";
			elsif QstateRE(2) = to_sfixed(02.1250,QstateRE(2)) then
				char2RE <= "+02.1250";
			elsif QstateRE(2) = to_sfixed(02.1875,QstateRE(2)) then
				char2RE <= "+02.1875";
			elsif QstateRE(2) = to_sfixed(02.2500,QstateRE(2)) then
				char2RE <= "+02.2500";
			elsif QstateRE(2) = to_sfixed(02.3125,QstateRE(2)) then
				char2RE <= "+02.3125";
			elsif QstateRE(2) = to_sfixed(02.3750,QstateRE(2)) then
				char2RE <= "+02.3750";
			elsif QstateRE(2) = to_sfixed(02.4375,QstateRE(2)) then
				char2RE <= "+02.4375";
			elsif QstateRE(2) = to_sfixed(02.5000,QstateRE(2)) then
				char2RE <= "+02.5000";
			elsif QstateRE(2) = to_sfixed(02.5625,QstateRE(2)) then
				char2RE <= "+02.5625";
			elsif QstateRE(2) = to_sfixed(02.6250,QstateRE(2)) then
				char2RE <= "+02.6250";
			elsif QstateRE(2) = to_sfixed(02.6875,QstateRE(2)) then
				char2RE <= "+02.6875";
			elsif QstateRE(2) = to_sfixed(02.7500,QstateRE(2)) then
				char2RE <= "+02.7500";
			elsif QstateRE(2) = to_sfixed(02.8125,QstateRE(2)) then
				char2RE <= "+02.8125";
			elsif QstateRE(2) = to_sfixed(02.8750,QstateRE(2)) then
				char2RE <= "+02.8750";
			elsif QstateRE(2) = to_sfixed(02.9375,QstateRE(2)) then
				char2RE <= "+02.9375";
			elsif QstateRE(2) = to_sfixed(03.0000,QstateRE(2)) then
				char2RE <= "+03.0000";
			elsif QstateRE(2) = to_sfixed(03.0625,QstateRE(2)) then
				char2RE <= "+03.0625";
			elsif QstateRE(2) = to_sfixed(03.1250,QstateRE(2)) then
				char2RE <= "+03.1250";
			elsif QstateRE(2) = to_sfixed(03.1875,QstateRE(2)) then
				char2RE <= "+03.1875";
			elsif QstateRE(2) = to_sfixed(03.2500,QstateRE(2)) then
				char2RE <= "+03.2500";
			elsif QstateRE(2) = to_sfixed(03.3125,QstateRE(2)) then
				char2RE <= "+03.3125";
			elsif QstateRE(2) = to_sfixed(03.3750,QstateRE(2)) then
				char2RE <= "+03.3750";
			elsif QstateRE(2) = to_sfixed(03.4375,QstateRE(2)) then
				char2RE <= "+03.4375";
			elsif QstateRE(2) = to_sfixed(03.5000,QstateRE(2)) then
				char2RE <= "+03.5000";
			elsif QstateRE(2) = to_sfixed(03.5625,QstateRE(2)) then
				char2RE <= "+03.5625";
			elsif QstateRE(2) = to_sfixed(03.6250,QstateRE(2)) then
				char2RE <= "+03.6250";
			elsif QstateRE(2) = to_sfixed(03.6875,QstateRE(2)) then
				char2RE <= "+03.6875";
			elsif QstateRE(2) = to_sfixed(03.7500,QstateRE(2)) then
				char2RE <= "+03.7500";
			elsif QstateRE(2) = to_sfixed(03.8125,QstateRE(2)) then
				char2RE <= "+03.8125";
			elsif QstateRE(2) = to_sfixed(03.8750,QstateRE(2)) then
				char2RE <= "+03.8750";
			elsif QstateRE(2) = to_sfixed(03.9375,QstateRE(2)) then
				char2RE <= "+03.9375";
			elsif QstateRE(2) = to_sfixed(04.0000,QstateRE(2)) then
				char2RE <= "+04.0000";
			elsif QstateRE(2) = to_sfixed(04.0625,QstateRE(2)) then
				char2RE <= "+04.0625";
			elsif QstateRE(2) = to_sfixed(04.1250,QstateRE(2)) then
				char2RE <= "+04.1250";
			elsif QstateRE(2) = to_sfixed(04.1875,QstateRE(2)) then
				char2RE <= "+04.1875";
			elsif QstateRE(2) = to_sfixed(04.2500,QstateRE(2)) then
				char2RE <= "+04.2500";
			elsif QstateRE(2) = to_sfixed(04.3125,QstateRE(2)) then
				char2RE <= "+04.3125";
			elsif QstateRE(2) = to_sfixed(04.3750,QstateRE(2)) then
				char2RE <= "+04.3750";
			elsif QstateRE(2) = to_sfixed(04.4375,QstateRE(2)) then
				char2RE <= "+04.4375";
			elsif QstateRE(2) = to_sfixed(04.5000,QstateRE(2)) then
				char2RE <= "+04.5000";
			elsif QstateRE(2) = to_sfixed(04.5625,QstateRE(2)) then
				char2RE <= "+04.5625";
			elsif QstateRE(2) = to_sfixed(04.6250,QstateRE(2)) then
				char2RE <= "+04.6250";
			elsif QstateRE(2) = to_sfixed(04.6875,QstateRE(2)) then
				char2RE <= "+04.6875";
			elsif QstateRE(2) = to_sfixed(04.7500,QstateRE(2)) then
				char2RE <= "+04.7500";
			elsif QstateRE(2) = to_sfixed(04.8125,QstateRE(2)) then
				char2RE <= "+04.8125";
			elsif QstateRE(2) = to_sfixed(04.8750,QstateRE(2)) then
				char2RE <= "+04.8750";
			elsif QstateRE(2) = to_sfixed(04.9375,QstateRE(2)) then
				char2RE <= "+04.9375";
			elsif QstateRE(2) = to_sfixed(05.0000,QstateRE(2)) then
				char2RE <= "+05.0000";
			elsif QstateRE(2) = to_sfixed(05.0625,QstateRE(2)) then
				char2RE <= "+05.0625";
			elsif QstateRE(2) = to_sfixed(05.1250,QstateRE(2)) then
				char2RE <= "+05.1250";
			elsif QstateRE(2) = to_sfixed(05.1875,QstateRE(2)) then
				char2RE <= "+05.1875";
			elsif QstateRE(2) = to_sfixed(05.2500,QstateRE(2)) then
				char2RE <= "+05.2500";
			elsif QstateRE(2) = to_sfixed(05.3125,QstateRE(2)) then
				char2RE <= "+05.3125";
			elsif QstateRE(2) = to_sfixed(05.3750,QstateRE(2)) then
				char2RE <= "+05.3750";
			elsif QstateRE(2) = to_sfixed(05.4375,QstateRE(2)) then
				char2RE <= "+05.4375";
			elsif QstateRE(2) = to_sfixed(05.5000,QstateRE(2)) then
				char2RE <= "+05.5000";
			elsif QstateRE(2) = to_sfixed(05.5625,QstateRE(2)) then
				char2RE <= "+05.5625";
			elsif QstateRE(2) = to_sfixed(05.6250,QstateRE(2)) then
				char2RE <= "+05.6250";
			elsif QstateRE(2) = to_sfixed(05.6875,QstateRE(2)) then
				char2RE <= "+05.6875";
			elsif QstateRE(2) = to_sfixed(05.7500,QstateRE(2)) then
				char2RE <= "+05.7500";
			elsif QstateRE(2) = to_sfixed(05.8125,QstateRE(2)) then
				char2RE <= "+05.8125";
			elsif QstateRE(2) = to_sfixed(05.8750,QstateRE(2)) then
				char2RE <= "+05.8750";
			elsif QstateRE(2) = to_sfixed(05.9375,QstateRE(2)) then
				char2RE <= "+05.9375";
			elsif QstateRE(2) = to_sfixed(06.0000,QstateRE(2)) then
				char2RE <= "+06.0000";
			elsif QstateRE(2) = to_sfixed(06.0625,QstateRE(2)) then
				char2RE <= "+06.0625";
			elsif QstateRE(2) = to_sfixed(06.1250,QstateRE(2)) then
				char2RE <= "+06.1250";
			elsif QstateRE(2) = to_sfixed(06.1875,QstateRE(2)) then
				char2RE <= "+06.1875";
			elsif QstateRE(2) = to_sfixed(06.2500,QstateRE(2)) then
				char2RE <= "+06.2500";
			elsif QstateRE(2) = to_sfixed(06.3125,QstateRE(2)) then
				char2RE <= "+06.3125";
			elsif QstateRE(2) = to_sfixed(06.3750,QstateRE(2)) then
				char2RE <= "+06.3750";
			elsif QstateRE(2) = to_sfixed(06.4375,QstateRE(2)) then
				char2RE <= "+06.4375";
			elsif QstateRE(2) = to_sfixed(06.5000,QstateRE(2)) then
				char2RE <= "+06.5000";
			elsif QstateRE(2) = to_sfixed(06.5625,QstateRE(2)) then
				char2RE <= "+06.5625";
			elsif QstateRE(2) = to_sfixed(06.6250,QstateRE(2)) then
				char2RE <= "+06.6250";
			elsif QstateRE(2) = to_sfixed(06.6875,QstateRE(2)) then
				char2RE <= "+06.6875";
			elsif QstateRE(2) = to_sfixed(06.7500,QstateRE(2)) then
				char2RE <= "+06.7500";
			elsif QstateRE(2) = to_sfixed(06.8125,QstateRE(2)) then
				char2RE <= "+06.8125";
			elsif QstateRE(2) = to_sfixed(06.8750,QstateRE(2)) then
				char2RE <= "+06.8750";
			elsif QstateRE(2) = to_sfixed(06.9375,QstateRE(2)) then
				char2RE <= "+06.9375";
			elsif QstateRE(2) = to_sfixed(07.0000,QstateRE(2)) then
				char2RE <= "+07.0000";
			elsif QstateRE(2) = to_sfixed(07.0625,QstateRE(2)) then
				char2RE <= "+07.0625";
			elsif QstateRE(2) = to_sfixed(07.1250,QstateRE(2)) then
				char2RE <= "+07.1250";
			elsif QstateRE(2) = to_sfixed(07.1875,QstateRE(2)) then
				char2RE <= "+07.1875";
			elsif QstateRE(2) = to_sfixed(07.2500,QstateRE(2)) then
				char2RE <= "+07.2500";
			elsif QstateRE(2) = to_sfixed(07.3125,QstateRE(2)) then
				char2RE <= "+07.3125";
			elsif QstateRE(2) = to_sfixed(07.3750,QstateRE(2)) then
				char2RE <= "+07.3750";
			elsif QstateRE(2) = to_sfixed(07.4375,QstateRE(2)) then
				char2RE <= "+07.4375";
			elsif QstateRE(2) = to_sfixed(07.5000,QstateRE(2)) then
				char2RE <= "+07.5000";
			elsif QstateRE(2) = to_sfixed(07.5625,QstateRE(2)) then
				char2RE <= "+07.5625";
			elsif QstateRE(2) = to_sfixed(07.6250,QstateRE(2)) then
				char2RE <= "+07.6250";
			elsif QstateRE(2) = to_sfixed(07.6875,QstateRE(2)) then
				char2RE <= "+07.6875";
			elsif QstateRE(2) = to_sfixed(07.7500,QstateRE(2)) then
				char2RE <= "+07.7500";
			elsif QstateRE(2) = to_sfixed(07.8125,QstateRE(2)) then
				char2RE <= "+07.8125";
			elsif QstateRE(2) = to_sfixed(07.8750,QstateRE(2)) then
				char2RE <= "+07.8750";
			elsif QstateRE(2) = to_sfixed(07.9375,QstateRE(2)) then
				char2RE <= "+07.9375";
			elsif QstateRE(2) = to_sfixed(08.0000,QstateRE(2)) then
				char2RE <= "+08.0000";
			elsif QstateRE(2) = to_sfixed(08.0625,QstateRE(2)) then
				char2RE <= "+08.0625";
			elsif QstateRE(2) = to_sfixed(08.1250,QstateRE(2)) then
				char2RE <= "+08.1250";
			elsif QstateRE(2) = to_sfixed(08.1875,QstateRE(2)) then
				char2RE <= "+08.1875";
			elsif QstateRE(2) = to_sfixed(08.2500,QstateRE(2)) then
				char2RE <= "+08.2500";
			elsif QstateRE(2) = to_sfixed(08.3125,QstateRE(2)) then
				char2RE <= "+08.3125";
			elsif QstateRE(2) = to_sfixed(08.3750,QstateRE(2)) then
				char2RE <= "+08.3750";
			elsif QstateRE(2) = to_sfixed(08.4375,QstateRE(2)) then
				char2RE <= "+08.4375";
			elsif QstateRE(2) = to_sfixed(08.5000,QstateRE(2)) then
				char2RE <= "+08.5000";
			elsif QstateRE(2) = to_sfixed(08.5625,QstateRE(2)) then
				char2RE <= "+08.5625";
			elsif QstateRE(2) = to_sfixed(08.6250,QstateRE(2)) then
				char2RE <= "+08.6250";
			elsif QstateRE(2) = to_sfixed(08.6875,QstateRE(2)) then
				char2RE <= "+08.6875";
			elsif QstateRE(2) = to_sfixed(08.7500,QstateRE(2)) then
				char2RE <= "+08.7500";
			elsif QstateRE(2) = to_sfixed(08.8125,QstateRE(2)) then
				char2RE <= "+08.8125";
			elsif QstateRE(2) = to_sfixed(08.8750,QstateRE(2)) then
				char2RE <= "+08.8750";
			elsif QstateRE(2) = to_sfixed(08.9375,QstateRE(2)) then
				char2RE <= "+08.9375";
			elsif QstateRE(2) = to_sfixed(09.0000,QstateRE(2)) then
				char2RE <= "+09.0000";
			elsif QstateRE(2) = to_sfixed(09.0625,QstateRE(2)) then
				char2RE <= "+09.0625";
			elsif QstateRE(2) = to_sfixed(09.1250,QstateRE(2)) then
				char2RE <= "+09.1250";
			elsif QstateRE(2) = to_sfixed(09.1875,QstateRE(2)) then
				char2RE <= "+09.1875";
			elsif QstateRE(2) = to_sfixed(09.2500,QstateRE(2)) then
				char2RE <= "+09.2500";
			elsif QstateRE(2) = to_sfixed(09.3125,QstateRE(2)) then
				char2RE <= "+09.3125";
			elsif QstateRE(2) = to_sfixed(09.3750,QstateRE(2)) then
				char2RE <= "+09.3750";
			elsif QstateRE(2) = to_sfixed(09.4375,QstateRE(2)) then
				char2RE <= "+09.4375";
			elsif QstateRE(2) = to_sfixed(09.5000,QstateRE(2)) then
				char2RE <= "+09.5000";
			elsif QstateRE(2) = to_sfixed(09.5625,QstateRE(2)) then
				char2RE <= "+09.5625";
			elsif QstateRE(2) = to_sfixed(09.6250,QstateRE(2)) then
				char2RE <= "+09.6250";
			elsif QstateRE(2) = to_sfixed(09.6875,QstateRE(2)) then
				char2RE <= "+09.6875";
			elsif QstateRE(2) = to_sfixed(09.7500,QstateRE(2)) then
				char2RE <= "+09.7500";
			elsif QstateRE(2) = to_sfixed(09.8125,QstateRE(2)) then
				char2RE <= "+09.8125";
			elsif QstateRE(2) = to_sfixed(09.8750,QstateRE(2)) then
				char2RE <= "+09.8750";
			elsif QstateRE(2) = to_sfixed(09.9375,QstateRE(2)) then
				char2RE <= "+09.9375";
			elsif QstateRE(2) = to_sfixed(10.0000,QstateRE(2)) then
				char2RE <= "+10.0000";
			elsif QstateRE(2) = to_sfixed(10.0625,QstateRE(2)) then
				char2RE <= "+10.0625";
			elsif QstateRE(2) = to_sfixed(10.1250,QstateRE(2)) then
				char2RE <= "+10.1250";
			elsif QstateRE(2) = to_sfixed(10.1875,QstateRE(2)) then
				char2RE <= "+10.1875";
			elsif QstateRE(2) = to_sfixed(10.2500,QstateRE(2)) then
				char2RE <= "+10.2500";
			elsif QstateRE(2) = to_sfixed(10.3125,QstateRE(2)) then
				char2RE <= "+10.3125";
			elsif QstateRE(2) = to_sfixed(10.3750,QstateRE(2)) then
				char2RE <= "+10.3750";
			elsif QstateRE(2) = to_sfixed(10.4375,QstateRE(2)) then
				char2RE <= "+10.4375";
			elsif QstateRE(2) = to_sfixed(10.5000,QstateRE(2)) then
				char2RE <= "+10.5000";
			elsif QstateRE(2) = to_sfixed(10.5625,QstateRE(2)) then
				char2RE <= "+10.5625";
			elsif QstateRE(2) = to_sfixed(10.6250,QstateRE(2)) then
				char2RE <= "+10.6250";
			elsif QstateRE(2) = to_sfixed(10.6875,QstateRE(2)) then
				char2RE <= "+10.6875";
			elsif QstateRE(2) = to_sfixed(10.7500,QstateRE(2)) then
				char2RE <= "+10.7500";
			elsif QstateRE(2) = to_sfixed(10.8125,QstateRE(2)) then
				char2RE <= "+10.8125";
			elsif QstateRE(2) = to_sfixed(10.8750,QstateRE(2)) then
				char2RE <= "+10.8750";
			elsif QstateRE(2) = to_sfixed(10.9375,QstateRE(2)) then
				char2RE <= "+10.9375";
			elsif QstateRE(2) = to_sfixed(11.0000,QstateRE(2)) then
				char2RE <= "+11.0000";
			elsif QstateRE(2) = to_sfixed(11.0625,QstateRE(2)) then
				char2RE <= "+11.0625";
			elsif QstateRE(2) = to_sfixed(11.1250,QstateRE(2)) then
				char2RE <= "+11.1250";
			elsif QstateRE(2) = to_sfixed(11.1875,QstateRE(2)) then
				char2RE <= "+11.1875";
			elsif QstateRE(2) = to_sfixed(11.2500,QstateRE(2)) then
				char2RE <= "+11.2500";
			elsif QstateRE(2) = to_sfixed(11.3125,QstateRE(2)) then
				char2RE <= "+11.3125";
			elsif QstateRE(2) = to_sfixed(11.3750,QstateRE(2)) then
				char2RE <= "+11.3750";
			elsif QstateRE(2) = to_sfixed(11.4375,QstateRE(2)) then
				char2RE <= "+11.4375";
			elsif QstateRE(2) = to_sfixed(11.5000,QstateRE(2)) then
				char2RE <= "+11.5000";
			elsif QstateRE(2) = to_sfixed(11.5625,QstateRE(2)) then
				char2RE <= "+11.5625";
			elsif QstateRE(2) = to_sfixed(11.6250,QstateRE(2)) then
				char2RE <= "+11.6250";
			elsif QstateRE(2) = to_sfixed(11.6875,QstateRE(2)) then
				char2RE <= "+11.6875";
			elsif QstateRE(2) = to_sfixed(11.7500,QstateRE(2)) then
				char2RE <= "+11.7500";
			elsif QstateRE(2) = to_sfixed(11.8125,QstateRE(2)) then
				char2RE <= "+11.8125";
			elsif QstateRE(2) = to_sfixed(11.8750,QstateRE(2)) then
				char2RE <= "+11.8750";
			elsif QstateRE(2) = to_sfixed(11.9375,QstateRE(2)) then
				char2RE <= "+11.9375";
			elsif QstateRE(2) = to_sfixed(12.0000,QstateRE(2)) then
				char2RE <= "+12.0000";
			elsif QstateRE(2) = to_sfixed(12.0625,QstateRE(2)) then
				char2RE <= "+12.0625";
			elsif QstateRE(2) = to_sfixed(12.1250,QstateRE(2)) then
				char2RE <= "+12.1250";
			elsif QstateRE(2) = to_sfixed(12.1875,QstateRE(2)) then
				char2RE <= "+12.1875";
			elsif QstateRE(2) = to_sfixed(12.2500,QstateRE(2)) then
				char2RE <= "+12.2500";
			elsif QstateRE(2) = to_sfixed(12.3125,QstateRE(2)) then
				char2RE <= "+12.3125";
			elsif QstateRE(2) = to_sfixed(12.3750,QstateRE(2)) then
				char2RE <= "+12.3750";
			elsif QstateRE(2) = to_sfixed(12.4375,QstateRE(2)) then
				char2RE <= "+12.4375";
			elsif QstateRE(2) = to_sfixed(12.5000,QstateRE(2)) then
				char2RE <= "+12.5000";
			elsif QstateRE(2) = to_sfixed(12.5625,QstateRE(2)) then
				char2RE <= "+12.5625";
			elsif QstateRE(2) = to_sfixed(12.6250,QstateRE(2)) then
				char2RE <= "+12.6250";
			elsif QstateRE(2) = to_sfixed(12.6875,QstateRE(2)) then
				char2RE <= "+12.6875";
			elsif QstateRE(2) = to_sfixed(12.7500,QstateRE(2)) then
				char2RE <= "+12.7500";
			elsif QstateRE(2) = to_sfixed(12.8125,QstateRE(2)) then
				char2RE <= "+12.8125";
			elsif QstateRE(2) = to_sfixed(12.8750,QstateRE(2)) then
				char2RE <= "+12.8750";
			elsif QstateRE(2) = to_sfixed(12.9375,QstateRE(2)) then
				char2RE <= "+12.9375";
			elsif QstateRE(2) = to_sfixed(13.0000,QstateRE(2)) then
				char2RE <= "+13.0000";
			elsif QstateRE(2) = to_sfixed(13.0625,QstateRE(2)) then
				char2RE <= "+13.0625";
			elsif QstateRE(2) = to_sfixed(13.1250,QstateRE(2)) then
				char2RE <= "+13.1250";
			elsif QstateRE(2) = to_sfixed(13.1875,QstateRE(2)) then
				char2RE <= "+13.1875";
			elsif QstateRE(2) = to_sfixed(13.2500,QstateRE(2)) then
				char2RE <= "+13.2500";
			elsif QstateRE(2) = to_sfixed(13.3125,QstateRE(2)) then
				char2RE <= "+13.3125";
			elsif QstateRE(2) = to_sfixed(13.3750,QstateRE(2)) then
				char2RE <= "+13.3750";
			elsif QstateRE(2) = to_sfixed(13.4375,QstateRE(2)) then
				char2RE <= "+13.4375";
			elsif QstateRE(2) = to_sfixed(13.5000,QstateRE(2)) then
				char2RE <= "+13.5000";
			elsif QstateRE(2) = to_sfixed(13.5625,QstateRE(2)) then
				char2RE <= "+13.5625";
			elsif QstateRE(2) = to_sfixed(13.6250,QstateRE(2)) then
				char2RE <= "+13.6250";
			elsif QstateRE(2) = to_sfixed(13.6875,QstateRE(2)) then
				char2RE <= "+13.6875";
			elsif QstateRE(2) = to_sfixed(13.7500,QstateRE(2)) then
				char2RE <= "+13.7500";
			elsif QstateRE(2) = to_sfixed(13.8125,QstateRE(2)) then
				char2RE <= "+13.8125";
			elsif QstateRE(2) = to_sfixed(13.8750,QstateRE(2)) then
				char2RE <= "+13.8750";
			elsif QstateRE(2) = to_sfixed(13.9375,QstateRE(2)) then
				char2RE <= "+13.9375";
			elsif QstateRE(2) = to_sfixed(14.0000,QstateRE(2)) then
				char2RE <= "+14.0000";
			elsif QstateRE(2) = to_sfixed(14.0625,QstateRE(2)) then
				char2RE <= "+14.0625";
			elsif QstateRE(2) = to_sfixed(14.1250,QstateRE(2)) then
				char2RE <= "+14.1250";
			elsif QstateRE(2) = to_sfixed(14.1875,QstateRE(2)) then
				char2RE <= "+14.1875";
			elsif QstateRE(2) = to_sfixed(14.2500,QstateRE(2)) then
				char2RE <= "+14.2500";
			elsif QstateRE(2) = to_sfixed(14.3125,QstateRE(2)) then
				char2RE <= "+14.3125";
			elsif QstateRE(2) = to_sfixed(14.3750,QstateRE(2)) then
				char2RE <= "+14.3750";
			elsif QstateRE(2) = to_sfixed(14.4375,QstateRE(2)) then
				char2RE <= "+14.4375";
			elsif QstateRE(2) = to_sfixed(14.5000,QstateRE(2)) then
				char2RE <= "+14.5000";
			elsif QstateRE(2) = to_sfixed(14.5625,QstateRE(2)) then
				char2RE <= "+14.5625";
			elsif QstateRE(2) = to_sfixed(14.6250,QstateRE(2)) then
				char2RE <= "+14.6250";
			elsif QstateRE(2) = to_sfixed(14.6875,QstateRE(2)) then
				char2RE <= "+14.6875";
			elsif QstateRE(2) = to_sfixed(14.7500,QstateRE(2)) then
				char2RE <= "+14.7500";
			elsif QstateRE(2) = to_sfixed(14.8125,QstateRE(2)) then
				char2RE <= "+14.8125";
			elsif QstateRE(2) = to_sfixed(14.8750,QstateRE(2)) then
				char2RE <= "+14.8750";
			elsif QstateRE(2) = to_sfixed(14.9375,QstateRE(2)) then
				char2RE <= "+14.9375";
			elsif QstateRE(2) = to_sfixed(15.0000,QstateRE(2)) then
				char2RE <= "+15.0000";
			elsif QstateRE(2) = to_sfixed(15.0625,QstateRE(2)) then
				char2RE <= "+15.0625";
			elsif QstateRE(2) = to_sfixed(15.1250,QstateRE(2)) then
				char2RE <= "+15.1250";
			elsif QstateRE(2) = to_sfixed(15.1875,QstateRE(2)) then
				char2RE <= "+15.1875";
			elsif QstateRE(2) = to_sfixed(15.2500,QstateRE(2)) then
				char2RE <= "+15.2500";
			elsif QstateRE(2) = to_sfixed(15.3125,QstateRE(2)) then
				char2RE <= "+15.3125";
			elsif QstateRE(2) = to_sfixed(15.3750,QstateRE(2)) then
				char2RE <= "+15.3750";
			elsif QstateRE(2) = to_sfixed(15.4375,QstateRE(2)) then
				char2RE <= "+15.4375";
			elsif QstateRE(2) = to_sfixed(15.5000,QstateRE(2)) then
				char2RE <= "+15.5000";
			elsif QstateRE(2) = to_sfixed(15.5625,QstateRE(2)) then
				char2RE <= "+15.5625";
			elsif QstateRE(2) = to_sfixed(15.6250,QstateRE(2)) then
				char2RE <= "+15.6250";
			elsif QstateRE(2) = to_sfixed(15.6875,QstateRE(2)) then
				char2RE <= "+15.6875";
			elsif QstateRE(2) = to_sfixed(15.7500,QstateRE(2)) then
				char2RE <= "+15.7500";
			elsif QstateRE(2) = to_sfixed(15.8125,QstateRE(2)) then
				char2RE <= "+15.8125";
			elsif QstateRE(2) = to_sfixed(15.8750,QstateRE(2)) then
				char2RE <= "+15.8750";
			elsif QstateRE(2) = to_sfixed(15.9375,QstateRE(2)) then
				char2RE <= "+15.9375";
			end if;
			if QstateIM(2) = to_sfixed(-15.9375,QstateIM(2)) then
				char2IM <= "-15.9375";
			elsif QstateIM(2) = to_sfixed(-15.8750,QstateIM(2)) then
				char2IM <= "-15.8750";
			elsif QstateIM(2) = to_sfixed(-15.8125,QstateIM(2)) then
				char2IM <= "-15.8125";
			elsif QstateIM(2) = to_sfixed(-15.7500,QstateIM(2)) then
				char2IM <= "-15.7500";
			elsif QstateIM(2) = to_sfixed(-15.6875,QstateIM(2)) then
				char2IM <= "-15.6875";
			elsif QstateIM(2) = to_sfixed(-15.6250,QstateIM(2)) then
				char2IM <= "-15.6250";
			elsif QstateIM(2) = to_sfixed(-15.5625,QstateIM(2)) then
				char2IM <= "-15.5625";
			elsif QstateIM(2) = to_sfixed(-15.5000,QstateIM(2)) then
				char2IM <= "-15.5000";
			elsif QstateIM(2) = to_sfixed(-15.4375,QstateIM(2)) then
				char2IM <= "-15.4375";
			elsif QstateIM(2) = to_sfixed(-15.3750,QstateIM(2)) then
				char2IM <= "-15.3750";
			elsif QstateIM(2) = to_sfixed(-15.3125,QstateIM(2)) then
				char2IM <= "-15.3125";
			elsif QstateIM(2) = to_sfixed(-15.2500,QstateIM(2)) then
				char2IM <= "-15.2500";
			elsif QstateIM(2) = to_sfixed(-15.1875,QstateIM(2)) then
				char2IM <= "-15.1875";
			elsif QstateIM(2) = to_sfixed(-15.1250,QstateIM(2)) then
				char2IM <= "-15.1250";
			elsif QstateIM(2) = to_sfixed(-15.0625,QstateIM(2)) then
				char2IM <= "-15.0625";
			elsif QstateIM(2) = to_sfixed(-15.0000,QstateIM(2)) then
				char2IM <= "-15.0000";
			elsif QstateIM(2) = to_sfixed(-14.9375,QstateIM(2)) then
				char2IM <= "-14.9375";
			elsif QstateIM(2) = to_sfixed(-14.8750,QstateIM(2)) then
				char2IM <= "-14.8750";
			elsif QstateIM(2) = to_sfixed(-14.8125,QstateIM(2)) then
				char2IM <= "-14.8125";
			elsif QstateIM(2) = to_sfixed(-14.7500,QstateIM(2)) then
				char2IM <= "-14.7500";
			elsif QstateIM(2) = to_sfixed(-14.6875,QstateIM(2)) then
				char2IM <= "-14.6875";
			elsif QstateIM(2) = to_sfixed(-14.6250,QstateIM(2)) then
				char2IM <= "-14.6250";
			elsif QstateIM(2) = to_sfixed(-14.5625,QstateIM(2)) then
				char2IM <= "-14.5625";
			elsif QstateIM(2) = to_sfixed(-14.5000,QstateIM(2)) then
				char2IM <= "-14.5000";
			elsif QstateIM(2) = to_sfixed(-14.4375,QstateIM(2)) then
				char2IM <= "-14.4375";
			elsif QstateIM(2) = to_sfixed(-14.3750,QstateIM(2)) then
				char2IM <= "-14.3750";
			elsif QstateIM(2) = to_sfixed(-14.3125,QstateIM(2)) then
				char2IM <= "-14.3125";
			elsif QstateIM(2) = to_sfixed(-14.2500,QstateIM(2)) then
				char2IM <= "-14.2500";
			elsif QstateIM(2) = to_sfixed(-14.1875,QstateIM(2)) then
				char2IM <= "-14.1875";
			elsif QstateIM(2) = to_sfixed(-14.1250,QstateIM(2)) then
				char2IM <= "-14.1250";
			elsif QstateIM(2) = to_sfixed(-14.0625,QstateIM(2)) then
				char2IM <= "-14.0625";
			elsif QstateIM(2) = to_sfixed(-14.0000,QstateIM(2)) then
				char2IM <= "-14.0000";
			elsif QstateIM(2) = to_sfixed(-13.9375,QstateIM(2)) then
				char2IM <= "-13.9375";
			elsif QstateIM(2) = to_sfixed(-13.8750,QstateIM(2)) then
				char2IM <= "-13.8750";
			elsif QstateIM(2) = to_sfixed(-13.8125,QstateIM(2)) then
				char2IM <= "-13.8125";
			elsif QstateIM(2) = to_sfixed(-13.7500,QstateIM(2)) then
				char2IM <= "-13.7500";
			elsif QstateIM(2) = to_sfixed(-13.6875,QstateIM(2)) then
				char2IM <= "-13.6875";
			elsif QstateIM(2) = to_sfixed(-13.6250,QstateIM(2)) then
				char2IM <= "-13.6250";
			elsif QstateIM(2) = to_sfixed(-13.5625,QstateIM(2)) then
				char2IM <= "-13.5625";
			elsif QstateIM(2) = to_sfixed(-13.5000,QstateIM(2)) then
				char2IM <= "-13.5000";
			elsif QstateIM(2) = to_sfixed(-13.4375,QstateIM(2)) then
				char2IM <= "-13.4375";
			elsif QstateIM(2) = to_sfixed(-13.3750,QstateIM(2)) then
				char2IM <= "-13.3750";
			elsif QstateIM(2) = to_sfixed(-13.3125,QstateIM(2)) then
				char2IM <= "-13.3125";
			elsif QstateIM(2) = to_sfixed(-13.2500,QstateIM(2)) then
				char2IM <= "-13.2500";
			elsif QstateIM(2) = to_sfixed(-13.1875,QstateIM(2)) then
				char2IM <= "-13.1875";
			elsif QstateIM(2) = to_sfixed(-13.1250,QstateIM(2)) then
				char2IM <= "-13.1250";
			elsif QstateIM(2) = to_sfixed(-13.0625,QstateIM(2)) then
				char2IM <= "-13.0625";
			elsif QstateIM(2) = to_sfixed(-13.0000,QstateIM(2)) then
				char2IM <= "-13.0000";
			elsif QstateIM(2) = to_sfixed(-12.9375,QstateIM(2)) then
				char2IM <= "-12.9375";
			elsif QstateIM(2) = to_sfixed(-12.8750,QstateIM(2)) then
				char2IM <= "-12.8750";
			elsif QstateIM(2) = to_sfixed(-12.8125,QstateIM(2)) then
				char2IM <= "-12.8125";
			elsif QstateIM(2) = to_sfixed(-12.7500,QstateIM(2)) then
				char2IM <= "-12.7500";
			elsif QstateIM(2) = to_sfixed(-12.6875,QstateIM(2)) then
				char2IM <= "-12.6875";
			elsif QstateIM(2) = to_sfixed(-12.6250,QstateIM(2)) then
				char2IM <= "-12.6250";
			elsif QstateIM(2) = to_sfixed(-12.5625,QstateIM(2)) then
				char2IM <= "-12.5625";
			elsif QstateIM(2) = to_sfixed(-12.5000,QstateIM(2)) then
				char2IM <= "-12.5000";
			elsif QstateIM(2) = to_sfixed(-12.4375,QstateIM(2)) then
				char2IM <= "-12.4375";
			elsif QstateIM(2) = to_sfixed(-12.3750,QstateIM(2)) then
				char2IM <= "-12.3750";
			elsif QstateIM(2) = to_sfixed(-12.3125,QstateIM(2)) then
				char2IM <= "-12.3125";
			elsif QstateIM(2) = to_sfixed(-12.2500,QstateIM(2)) then
				char2IM <= "-12.2500";
			elsif QstateIM(2) = to_sfixed(-12.1875,QstateIM(2)) then
				char2IM <= "-12.1875";
			elsif QstateIM(2) = to_sfixed(-12.1250,QstateIM(2)) then
				char2IM <= "-12.1250";
			elsif QstateIM(2) = to_sfixed(-12.0625,QstateIM(2)) then
				char2IM <= "-12.0625";
			elsif QstateIM(2) = to_sfixed(-12.0000,QstateIM(2)) then
				char2IM <= "-12.0000";
			elsif QstateIM(2) = to_sfixed(-11.9375,QstateIM(2)) then
				char2IM <= "-11.9375";
			elsif QstateIM(2) = to_sfixed(-11.8750,QstateIM(2)) then
				char2IM <= "-11.8750";
			elsif QstateIM(2) = to_sfixed(-11.8125,QstateIM(2)) then
				char2IM <= "-11.8125";
			elsif QstateIM(2) = to_sfixed(-11.7500,QstateIM(2)) then
				char2IM <= "-11.7500";
			elsif QstateIM(2) = to_sfixed(-11.6875,QstateIM(2)) then
				char2IM <= "-11.6875";
			elsif QstateIM(2) = to_sfixed(-11.6250,QstateIM(2)) then
				char2IM <= "-11.6250";
			elsif QstateIM(2) = to_sfixed(-11.5625,QstateIM(2)) then
				char2IM <= "-11.5625";
			elsif QstateIM(2) = to_sfixed(-11.5000,QstateIM(2)) then
				char2IM <= "-11.5000";
			elsif QstateIM(2) = to_sfixed(-11.4375,QstateIM(2)) then
				char2IM <= "-11.4375";
			elsif QstateIM(2) = to_sfixed(-11.3750,QstateIM(2)) then
				char2IM <= "-11.3750";
			elsif QstateIM(2) = to_sfixed(-11.3125,QstateIM(2)) then
				char2IM <= "-11.3125";
			elsif QstateIM(2) = to_sfixed(-11.2500,QstateIM(2)) then
				char2IM <= "-11.2500";
			elsif QstateIM(2) = to_sfixed(-11.1875,QstateIM(2)) then
				char2IM <= "-11.1875";
			elsif QstateIM(2) = to_sfixed(-11.1250,QstateIM(2)) then
				char2IM <= "-11.1250";
			elsif QstateIM(2) = to_sfixed(-11.0625,QstateIM(2)) then
				char2IM <= "-11.0625";
			elsif QstateIM(2) = to_sfixed(-11.0000,QstateIM(2)) then
				char2IM <= "-11.0000";
			elsif QstateIM(2) = to_sfixed(-10.9375,QstateIM(2)) then
				char2IM <= "-10.9375";
			elsif QstateIM(2) = to_sfixed(-10.8750,QstateIM(2)) then
				char2IM <= "-10.8750";
			elsif QstateIM(2) = to_sfixed(-10.8125,QstateIM(2)) then
				char2IM <= "-10.8125";
			elsif QstateIM(2) = to_sfixed(-10.7500,QstateIM(2)) then
				char2IM <= "-10.7500";
			elsif QstateIM(2) = to_sfixed(-10.6875,QstateIM(2)) then
				char2IM <= "-10.6875";
			elsif QstateIM(2) = to_sfixed(-10.6250,QstateIM(2)) then
				char2IM <= "-10.6250";
			elsif QstateIM(2) = to_sfixed(-10.5625,QstateIM(2)) then
				char2IM <= "-10.5625";
			elsif QstateIM(2) = to_sfixed(-10.5000,QstateIM(2)) then
				char2IM <= "-10.5000";
			elsif QstateIM(2) = to_sfixed(-10.4375,QstateIM(2)) then
				char2IM <= "-10.4375";
			elsif QstateIM(2) = to_sfixed(-10.3750,QstateIM(2)) then
				char2IM <= "-10.3750";
			elsif QstateIM(2) = to_sfixed(-10.3125,QstateIM(2)) then
				char2IM <= "-10.3125";
			elsif QstateIM(2) = to_sfixed(-10.2500,QstateIM(2)) then
				char2IM <= "-10.2500";
			elsif QstateIM(2) = to_sfixed(-10.1875,QstateIM(2)) then
				char2IM <= "-10.1875";
			elsif QstateIM(2) = to_sfixed(-10.1250,QstateIM(2)) then
				char2IM <= "-10.1250";
			elsif QstateIM(2) = to_sfixed(-10.0625,QstateIM(2)) then
				char2IM <= "-10.0625";
			elsif QstateIM(2) = to_sfixed(-10.0000,QstateIM(2)) then
				char2IM <= "-10.0000";
			elsif QstateIM(2) = to_sfixed(-9.9375,QstateIM(2)) then
				char2IM <= "--9.9375";
			elsif QstateIM(2) = to_sfixed(-9.8750,QstateIM(2)) then
				char2IM <= "--9.8750";
			elsif QstateIM(2) = to_sfixed(-9.8125,QstateIM(2)) then
				char2IM <= "--9.8125";
			elsif QstateIM(2) = to_sfixed(-9.7500,QstateIM(2)) then
				char2IM <= "--9.7500";
			elsif QstateIM(2) = to_sfixed(-9.6875,QstateIM(2)) then
				char2IM <= "--9.6875";
			elsif QstateIM(2) = to_sfixed(-9.6250,QstateIM(2)) then
				char2IM <= "--9.6250";
			elsif QstateIM(2) = to_sfixed(-9.5625,QstateIM(2)) then
				char2IM <= "--9.5625";
			elsif QstateIM(2) = to_sfixed(-9.5000,QstateIM(2)) then
				char2IM <= "--9.5000";
			elsif QstateIM(2) = to_sfixed(-9.4375,QstateIM(2)) then
				char2IM <= "--9.4375";
			elsif QstateIM(2) = to_sfixed(-9.3750,QstateIM(2)) then
				char2IM <= "--9.3750";
			elsif QstateIM(2) = to_sfixed(-9.3125,QstateIM(2)) then
				char2IM <= "--9.3125";
			elsif QstateIM(2) = to_sfixed(-9.2500,QstateIM(2)) then
				char2IM <= "--9.2500";
			elsif QstateIM(2) = to_sfixed(-9.1875,QstateIM(2)) then
				char2IM <= "--9.1875";
			elsif QstateIM(2) = to_sfixed(-9.1250,QstateIM(2)) then
				char2IM <= "--9.1250";
			elsif QstateIM(2) = to_sfixed(-9.0625,QstateIM(2)) then
				char2IM <= "--9.0625";
			elsif QstateIM(2) = to_sfixed(-9.0000,QstateIM(2)) then
				char2IM <= "--9.0000";
			elsif QstateIM(2) = to_sfixed(-8.9375,QstateIM(2)) then
				char2IM <= "--8.9375";
			elsif QstateIM(2) = to_sfixed(-8.8750,QstateIM(2)) then
				char2IM <= "--8.8750";
			elsif QstateIM(2) = to_sfixed(-8.8125,QstateIM(2)) then
				char2IM <= "--8.8125";
			elsif QstateIM(2) = to_sfixed(-8.7500,QstateIM(2)) then
				char2IM <= "--8.7500";
			elsif QstateIM(2) = to_sfixed(-8.6875,QstateIM(2)) then
				char2IM <= "--8.6875";
			elsif QstateIM(2) = to_sfixed(-8.6250,QstateIM(2)) then
				char2IM <= "--8.6250";
			elsif QstateIM(2) = to_sfixed(-8.5625,QstateIM(2)) then
				char2IM <= "--8.5625";
			elsif QstateIM(2) = to_sfixed(-8.5000,QstateIM(2)) then
				char2IM <= "--8.5000";
			elsif QstateIM(2) = to_sfixed(-8.4375,QstateIM(2)) then
				char2IM <= "--8.4375";
			elsif QstateIM(2) = to_sfixed(-8.3750,QstateIM(2)) then
				char2IM <= "--8.3750";
			elsif QstateIM(2) = to_sfixed(-8.3125,QstateIM(2)) then
				char2IM <= "--8.3125";
			elsif QstateIM(2) = to_sfixed(-8.2500,QstateIM(2)) then
				char2IM <= "--8.2500";
			elsif QstateIM(2) = to_sfixed(-8.1875,QstateIM(2)) then
				char2IM <= "--8.1875";
			elsif QstateIM(2) = to_sfixed(-8.1250,QstateIM(2)) then
				char2IM <= "--8.1250";
			elsif QstateIM(2) = to_sfixed(-8.0625,QstateIM(2)) then
				char2IM <= "--8.0625";
			elsif QstateIM(2) = to_sfixed(-8.0000,QstateIM(2)) then
				char2IM <= "--8.0000";
			elsif QstateIM(2) = to_sfixed(-7.9375,QstateIM(2)) then
				char2IM <= "--7.9375";
			elsif QstateIM(2) = to_sfixed(-7.8750,QstateIM(2)) then
				char2IM <= "--7.8750";
			elsif QstateIM(2) = to_sfixed(-7.8125,QstateIM(2)) then
				char2IM <= "--7.8125";
			elsif QstateIM(2) = to_sfixed(-7.7500,QstateIM(2)) then
				char2IM <= "--7.7500";
			elsif QstateIM(2) = to_sfixed(-7.6875,QstateIM(2)) then
				char2IM <= "--7.6875";
			elsif QstateIM(2) = to_sfixed(-7.6250,QstateIM(2)) then
				char2IM <= "--7.6250";
			elsif QstateIM(2) = to_sfixed(-7.5625,QstateIM(2)) then
				char2IM <= "--7.5625";
			elsif QstateIM(2) = to_sfixed(-7.5000,QstateIM(2)) then
				char2IM <= "--7.5000";
			elsif QstateIM(2) = to_sfixed(-7.4375,QstateIM(2)) then
				char2IM <= "--7.4375";
			elsif QstateIM(2) = to_sfixed(-7.3750,QstateIM(2)) then
				char2IM <= "--7.3750";
			elsif QstateIM(2) = to_sfixed(-7.3125,QstateIM(2)) then
				char2IM <= "--7.3125";
			elsif QstateIM(2) = to_sfixed(-7.2500,QstateIM(2)) then
				char2IM <= "--7.2500";
			elsif QstateIM(2) = to_sfixed(-7.1875,QstateIM(2)) then
				char2IM <= "--7.1875";
			elsif QstateIM(2) = to_sfixed(-7.1250,QstateIM(2)) then
				char2IM <= "--7.1250";
			elsif QstateIM(2) = to_sfixed(-7.0625,QstateIM(2)) then
				char2IM <= "--7.0625";
			elsif QstateIM(2) = to_sfixed(-7.0000,QstateIM(2)) then
				char2IM <= "--7.0000";
			elsif QstateIM(2) = to_sfixed(-6.9375,QstateIM(2)) then
				char2IM <= "--6.9375";
			elsif QstateIM(2) = to_sfixed(-6.8750,QstateIM(2)) then
				char2IM <= "--6.8750";
			elsif QstateIM(2) = to_sfixed(-6.8125,QstateIM(2)) then
				char2IM <= "--6.8125";
			elsif QstateIM(2) = to_sfixed(-6.7500,QstateIM(2)) then
				char2IM <= "--6.7500";
			elsif QstateIM(2) = to_sfixed(-6.6875,QstateIM(2)) then
				char2IM <= "--6.6875";
			elsif QstateIM(2) = to_sfixed(-6.6250,QstateIM(2)) then
				char2IM <= "--6.6250";
			elsif QstateIM(2) = to_sfixed(-6.5625,QstateIM(2)) then
				char2IM <= "--6.5625";
			elsif QstateIM(2) = to_sfixed(-6.5000,QstateIM(2)) then
				char2IM <= "--6.5000";
			elsif QstateIM(2) = to_sfixed(-6.4375,QstateIM(2)) then
				char2IM <= "--6.4375";
			elsif QstateIM(2) = to_sfixed(-6.3750,QstateIM(2)) then
				char2IM <= "--6.3750";
			elsif QstateIM(2) = to_sfixed(-6.3125,QstateIM(2)) then
				char2IM <= "--6.3125";
			elsif QstateIM(2) = to_sfixed(-6.2500,QstateIM(2)) then
				char2IM <= "--6.2500";
			elsif QstateIM(2) = to_sfixed(-6.1875,QstateIM(2)) then
				char2IM <= "--6.1875";
			elsif QstateIM(2) = to_sfixed(-6.1250,QstateIM(2)) then
				char2IM <= "--6.1250";
			elsif QstateIM(2) = to_sfixed(-6.0625,QstateIM(2)) then
				char2IM <= "--6.0625";
			elsif QstateIM(2) = to_sfixed(-6.0000,QstateIM(2)) then
				char2IM <= "--6.0000";
			elsif QstateIM(2) = to_sfixed(-5.9375,QstateIM(2)) then
				char2IM <= "--5.9375";
			elsif QstateIM(2) = to_sfixed(-5.8750,QstateIM(2)) then
				char2IM <= "--5.8750";
			elsif QstateIM(2) = to_sfixed(-5.8125,QstateIM(2)) then
				char2IM <= "--5.8125";
			elsif QstateIM(2) = to_sfixed(-5.7500,QstateIM(2)) then
				char2IM <= "--5.7500";
			elsif QstateIM(2) = to_sfixed(-5.6875,QstateIM(2)) then
				char2IM <= "--5.6875";
			elsif QstateIM(2) = to_sfixed(-5.6250,QstateIM(2)) then
				char2IM <= "--5.6250";
			elsif QstateIM(2) = to_sfixed(-5.5625,QstateIM(2)) then
				char2IM <= "--5.5625";
			elsif QstateIM(2) = to_sfixed(-5.5000,QstateIM(2)) then
				char2IM <= "--5.5000";
			elsif QstateIM(2) = to_sfixed(-5.4375,QstateIM(2)) then
				char2IM <= "--5.4375";
			elsif QstateIM(2) = to_sfixed(-5.3750,QstateIM(2)) then
				char2IM <= "--5.3750";
			elsif QstateIM(2) = to_sfixed(-5.3125,QstateIM(2)) then
				char2IM <= "--5.3125";
			elsif QstateIM(2) = to_sfixed(-5.2500,QstateIM(2)) then
				char2IM <= "--5.2500";
			elsif QstateIM(2) = to_sfixed(-5.1875,QstateIM(2)) then
				char2IM <= "--5.1875";
			elsif QstateIM(2) = to_sfixed(-5.1250,QstateIM(2)) then
				char2IM <= "--5.1250";
			elsif QstateIM(2) = to_sfixed(-5.0625,QstateIM(2)) then
				char2IM <= "--5.0625";
			elsif QstateIM(2) = to_sfixed(-5.0000,QstateIM(2)) then
				char2IM <= "--5.0000";
			elsif QstateIM(2) = to_sfixed(-4.9375,QstateIM(2)) then
				char2IM <= "--4.9375";
			elsif QstateIM(2) = to_sfixed(-4.8750,QstateIM(2)) then
				char2IM <= "--4.8750";
			elsif QstateIM(2) = to_sfixed(-4.8125,QstateIM(2)) then
				char2IM <= "--4.8125";
			elsif QstateIM(2) = to_sfixed(-4.7500,QstateIM(2)) then
				char2IM <= "--4.7500";
			elsif QstateIM(2) = to_sfixed(-4.6875,QstateIM(2)) then
				char2IM <= "--4.6875";
			elsif QstateIM(2) = to_sfixed(-4.6250,QstateIM(2)) then
				char2IM <= "--4.6250";
			elsif QstateIM(2) = to_sfixed(-4.5625,QstateIM(2)) then
				char2IM <= "--4.5625";
			elsif QstateIM(2) = to_sfixed(-4.5000,QstateIM(2)) then
				char2IM <= "--4.5000";
			elsif QstateIM(2) = to_sfixed(-4.4375,QstateIM(2)) then
				char2IM <= "--4.4375";
			elsif QstateIM(2) = to_sfixed(-4.3750,QstateIM(2)) then
				char2IM <= "--4.3750";
			elsif QstateIM(2) = to_sfixed(-4.3125,QstateIM(2)) then
				char2IM <= "--4.3125";
			elsif QstateIM(2) = to_sfixed(-4.2500,QstateIM(2)) then
				char2IM <= "--4.2500";
			elsif QstateIM(2) = to_sfixed(-4.1875,QstateIM(2)) then
				char2IM <= "--4.1875";
			elsif QstateIM(2) = to_sfixed(-4.1250,QstateIM(2)) then
				char2IM <= "--4.1250";
			elsif QstateIM(2) = to_sfixed(-4.0625,QstateIM(2)) then
				char2IM <= "--4.0625";
			elsif QstateIM(2) = to_sfixed(-4.0000,QstateIM(2)) then
				char2IM <= "--4.0000";
			elsif QstateIM(2) = to_sfixed(-3.9375,QstateIM(2)) then
				char2IM <= "--3.9375";
			elsif QstateIM(2) = to_sfixed(-3.8750,QstateIM(2)) then
				char2IM <= "--3.8750";
			elsif QstateIM(2) = to_sfixed(-3.8125,QstateIM(2)) then
				char2IM <= "--3.8125";
			elsif QstateIM(2) = to_sfixed(-3.7500,QstateIM(2)) then
				char2IM <= "--3.7500";
			elsif QstateIM(2) = to_sfixed(-3.6875,QstateIM(2)) then
				char2IM <= "--3.6875";
			elsif QstateIM(2) = to_sfixed(-3.6250,QstateIM(2)) then
				char2IM <= "--3.6250";
			elsif QstateIM(2) = to_sfixed(-3.5625,QstateIM(2)) then
				char2IM <= "--3.5625";
			elsif QstateIM(2) = to_sfixed(-3.5000,QstateIM(2)) then
				char2IM <= "--3.5000";
			elsif QstateIM(2) = to_sfixed(-3.4375,QstateIM(2)) then
				char2IM <= "--3.4375";
			elsif QstateIM(2) = to_sfixed(-3.3750,QstateIM(2)) then
				char2IM <= "--3.3750";
			elsif QstateIM(2) = to_sfixed(-3.3125,QstateIM(2)) then
				char2IM <= "--3.3125";
			elsif QstateIM(2) = to_sfixed(-3.2500,QstateIM(2)) then
				char2IM <= "--3.2500";
			elsif QstateIM(2) = to_sfixed(-3.1875,QstateIM(2)) then
				char2IM <= "--3.1875";
			elsif QstateIM(2) = to_sfixed(-3.1250,QstateIM(2)) then
				char2IM <= "--3.1250";
			elsif QstateIM(2) = to_sfixed(-3.0625,QstateIM(2)) then
				char2IM <= "--3.0625";
			elsif QstateIM(2) = to_sfixed(-3.0000,QstateIM(2)) then
				char2IM <= "--3.0000";
			elsif QstateIM(2) = to_sfixed(-2.9375,QstateIM(2)) then
				char2IM <= "--2.9375";
			elsif QstateIM(2) = to_sfixed(-2.8750,QstateIM(2)) then
				char2IM <= "--2.8750";
			elsif QstateIM(2) = to_sfixed(-2.8125,QstateIM(2)) then
				char2IM <= "--2.8125";
			elsif QstateIM(2) = to_sfixed(-2.7500,QstateIM(2)) then
				char2IM <= "--2.7500";
			elsif QstateIM(2) = to_sfixed(-2.6875,QstateIM(2)) then
				char2IM <= "--2.6875";
			elsif QstateIM(2) = to_sfixed(-2.6250,QstateIM(2)) then
				char2IM <= "--2.6250";
			elsif QstateIM(2) = to_sfixed(-2.5625,QstateIM(2)) then
				char2IM <= "--2.5625";
			elsif QstateIM(2) = to_sfixed(-2.5000,QstateIM(2)) then
				char2IM <= "--2.5000";
			elsif QstateIM(2) = to_sfixed(-2.4375,QstateIM(2)) then
				char2IM <= "--2.4375";
			elsif QstateIM(2) = to_sfixed(-2.3750,QstateIM(2)) then
				char2IM <= "--2.3750";
			elsif QstateIM(2) = to_sfixed(-2.3125,QstateIM(2)) then
				char2IM <= "--2.3125";
			elsif QstateIM(2) = to_sfixed(-2.2500,QstateIM(2)) then
				char2IM <= "--2.2500";
			elsif QstateIM(2) = to_sfixed(-2.1875,QstateIM(2)) then
				char2IM <= "--2.1875";
			elsif QstateIM(2) = to_sfixed(-2.1250,QstateIM(2)) then
				char2IM <= "--2.1250";
			elsif QstateIM(2) = to_sfixed(-2.0625,QstateIM(2)) then
				char2IM <= "--2.0625";
			elsif QstateIM(2) = to_sfixed(-2.0000,QstateIM(2)) then
				char2IM <= "--2.0000";
			elsif QstateIM(2) = to_sfixed(-1.9375,QstateIM(2)) then
				char2IM <= "--1.9375";
			elsif QstateIM(2) = to_sfixed(-1.8750,QstateIM(2)) then
				char2IM <= "--1.8750";
			elsif QstateIM(2) = to_sfixed(-1.8125,QstateIM(2)) then
				char2IM <= "--1.8125";
			elsif QstateIM(2) = to_sfixed(-1.7500,QstateIM(2)) then
				char2IM <= "--1.7500";
			elsif QstateIM(2) = to_sfixed(-1.6875,QstateIM(2)) then
				char2IM <= "--1.6875";
			elsif QstateIM(2) = to_sfixed(-1.6250,QstateIM(2)) then
				char2IM <= "--1.6250";
			elsif QstateIM(2) = to_sfixed(-1.5625,QstateIM(2)) then
				char2IM <= "--1.5625";
			elsif QstateIM(2) = to_sfixed(-1.5000,QstateIM(2)) then
				char2IM <= "--1.5000";
			elsif QstateIM(2) = to_sfixed(-1.4375,QstateIM(2)) then
				char2IM <= "--1.4375";
			elsif QstateIM(2) = to_sfixed(-1.3750,QstateIM(2)) then
				char2IM <= "--1.3750";
			elsif QstateIM(2) = to_sfixed(-1.3125,QstateIM(2)) then
				char2IM <= "--1.3125";
			elsif QstateIM(2) = to_sfixed(-1.2500,QstateIM(2)) then
				char2IM <= "--1.2500";
			elsif QstateIM(2) = to_sfixed(-1.1875,QstateIM(2)) then
				char2IM <= "--1.1875";
			elsif QstateIM(2) = to_sfixed(-1.1250,QstateIM(2)) then
				char2IM <= "--1.1250";
			elsif QstateIM(2) = to_sfixed(-1.0625,QstateIM(2)) then
				char2IM <= "--1.0625";
			elsif QstateIM(2) = to_sfixed(-1.0000,QstateIM(2)) then
				char2IM <= "--1.0000";
			elsif QstateIM(2) = to_sfixed(-0.9375,QstateIM(2)) then
				char2IM <= "--0.9375";
			elsif QstateIM(2) = to_sfixed(-0.8750,QstateIM(2)) then
				char2IM <= "--0.8750";
			elsif QstateIM(2) = to_sfixed(-0.8125,QstateIM(2)) then
				char2IM <= "--0.8125";
			elsif QstateIM(2) = to_sfixed(-0.7500,QstateIM(2)) then
				char2IM <= "--0.7500";
			elsif QstateIM(2) = to_sfixed(-0.6875,QstateIM(2)) then
				char2IM <= "--0.6875";
			elsif QstateIM(2) = to_sfixed(-0.6250,QstateIM(2)) then
				char2IM <= "--0.6250";
			elsif QstateIM(2) = to_sfixed(-0.5625,QstateIM(2)) then
				char2IM <= "--0.5625";
			elsif QstateIM(2) = to_sfixed(-0.5000,QstateIM(2)) then
				char2IM <= "--0.5000";
			elsif QstateIM(2) = to_sfixed(-0.4375,QstateIM(2)) then
				char2IM <= "--0.4375";
			elsif QstateIM(2) = to_sfixed(-0.3750,QstateIM(2)) then
				char2IM <= "--0.3750";
			elsif QstateIM(2) = to_sfixed(-0.3125,QstateIM(2)) then
				char2IM <= "--0.3125";
			elsif QstateIM(2) = to_sfixed(-0.2500,QstateIM(2)) then
				char2IM <= "--0.2500";
			elsif QstateIM(2) = to_sfixed(-0.1875,QstateIM(2)) then
				char2IM <= "--0.1875";
			elsif QstateIM(2) = to_sfixed(-0.1250,QstateIM(2)) then
				char2IM <= "--0.1250";
			elsif QstateIM(2) = to_sfixed(-0.0625,QstateIM(2)) then
				char2IM <= "--0.0625";
			elsif QstateIM(2) = to_sfixed(00.0000,QstateIM(2)) then
				char2IM <= "+00.0000";
			elsif QstateIM(2) = to_sfixed(00.0625,QstateIM(2)) then
				char2IM <= "+00.0625";
			elsif QstateIM(2) = to_sfixed(00.1250,QstateIM(2)) then
				char2IM <= "+00.1250";
			elsif QstateIM(2) = to_sfixed(00.1875,QstateIM(2)) then
				char2IM <= "+00.1875";
			elsif QstateIM(2) = to_sfixed(00.2500,QstateIM(2)) then
				char2IM <= "+00.2500";
			elsif QstateIM(2) = to_sfixed(00.3125,QstateIM(2)) then
				char2IM <= "+00.3125";
			elsif QstateIM(2) = to_sfixed(00.3750,QstateIM(2)) then
				char2IM <= "+00.3750";
			elsif QstateIM(2) = to_sfixed(00.4375,QstateIM(2)) then
				char2IM <= "+00.4375";
			elsif QstateIM(2) = to_sfixed(00.5000,QstateIM(2)) then
				char2IM <= "+00.5000";
			elsif QstateIM(2) = to_sfixed(00.5625,QstateIM(2)) then
				char2IM <= "+00.5625";
			elsif QstateIM(2) = to_sfixed(00.6250,QstateIM(2)) then
				char2IM <= "+00.6250";
			elsif QstateIM(2) = to_sfixed(00.6875,QstateIM(2)) then
				char2IM <= "+00.6875";
			elsif QstateIM(2) = to_sfixed(00.7500,QstateIM(2)) then
				char2IM <= "+00.7500";
			elsif QstateIM(2) = to_sfixed(00.8125,QstateIM(2)) then
				char2IM <= "+00.8125";
			elsif QstateIM(2) = to_sfixed(00.8750,QstateIM(2)) then
				char2IM <= "+00.8750";
			elsif QstateIM(2) = to_sfixed(00.9375,QstateIM(2)) then
				char2IM <= "+00.9375";
			elsif QstateIM(2) = to_sfixed(01.0000,QstateIM(2)) then
				char2IM <= "+01.0000";
			elsif QstateIM(2) = to_sfixed(01.0625,QstateIM(2)) then
				char2IM <= "+01.0625";
			elsif QstateIM(2) = to_sfixed(01.1250,QstateIM(2)) then
				char2IM <= "+01.1250";
			elsif QstateIM(2) = to_sfixed(01.1875,QstateIM(2)) then
				char2IM <= "+01.1875";
			elsif QstateIM(2) = to_sfixed(01.2500,QstateIM(2)) then
				char2IM <= "+01.2500";
			elsif QstateIM(2) = to_sfixed(01.3125,QstateIM(2)) then
				char2IM <= "+01.3125";
			elsif QstateIM(2) = to_sfixed(01.3750,QstateIM(2)) then
				char2IM <= "+01.3750";
			elsif QstateIM(2) = to_sfixed(01.4375,QstateIM(2)) then
				char2IM <= "+01.4375";
			elsif QstateIM(2) = to_sfixed(01.5000,QstateIM(2)) then
				char2IM <= "+01.5000";
			elsif QstateIM(2) = to_sfixed(01.5625,QstateIM(2)) then
				char2IM <= "+01.5625";
			elsif QstateIM(2) = to_sfixed(01.6250,QstateIM(2)) then
				char2IM <= "+01.6250";
			elsif QstateIM(2) = to_sfixed(01.6875,QstateIM(2)) then
				char2IM <= "+01.6875";
			elsif QstateIM(2) = to_sfixed(01.7500,QstateIM(2)) then
				char2IM <= "+01.7500";
			elsif QstateIM(2) = to_sfixed(01.8125,QstateIM(2)) then
				char2IM <= "+01.8125";
			elsif QstateIM(2) = to_sfixed(01.8750,QstateIM(2)) then
				char2IM <= "+01.8750";
			elsif QstateIM(2) = to_sfixed(01.9375,QstateIM(2)) then
				char2IM <= "+01.9375";
			elsif QstateIM(2) = to_sfixed(02.0000,QstateIM(2)) then
				char2IM <= "+02.0000";
			elsif QstateIM(2) = to_sfixed(02.0625,QstateIM(2)) then
				char2IM <= "+02.0625";
			elsif QstateIM(2) = to_sfixed(02.1250,QstateIM(2)) then
				char2IM <= "+02.1250";
			elsif QstateIM(2) = to_sfixed(02.1875,QstateIM(2)) then
				char2IM <= "+02.1875";
			elsif QstateIM(2) = to_sfixed(02.2500,QstateIM(2)) then
				char2IM <= "+02.2500";
			elsif QstateIM(2) = to_sfixed(02.3125,QstateIM(2)) then
				char2IM <= "+02.3125";
			elsif QstateIM(2) = to_sfixed(02.3750,QstateIM(2)) then
				char2IM <= "+02.3750";
			elsif QstateIM(2) = to_sfixed(02.4375,QstateIM(2)) then
				char2IM <= "+02.4375";
			elsif QstateIM(2) = to_sfixed(02.5000,QstateIM(2)) then
				char2IM <= "+02.5000";
			elsif QstateIM(2) = to_sfixed(02.5625,QstateIM(2)) then
				char2IM <= "+02.5625";
			elsif QstateIM(2) = to_sfixed(02.6250,QstateIM(2)) then
				char2IM <= "+02.6250";
			elsif QstateIM(2) = to_sfixed(02.6875,QstateIM(2)) then
				char2IM <= "+02.6875";
			elsif QstateIM(2) = to_sfixed(02.7500,QstateIM(2)) then
				char2IM <= "+02.7500";
			elsif QstateIM(2) = to_sfixed(02.8125,QstateIM(2)) then
				char2IM <= "+02.8125";
			elsif QstateIM(2) = to_sfixed(02.8750,QstateIM(2)) then
				char2IM <= "+02.8750";
			elsif QstateIM(2) = to_sfixed(02.9375,QstateIM(2)) then
				char2IM <= "+02.9375";
			elsif QstateIM(2) = to_sfixed(03.0000,QstateIM(2)) then
				char2IM <= "+03.0000";
			elsif QstateIM(2) = to_sfixed(03.0625,QstateIM(2)) then
				char2IM <= "+03.0625";
			elsif QstateIM(2) = to_sfixed(03.1250,QstateIM(2)) then
				char2IM <= "+03.1250";
			elsif QstateIM(2) = to_sfixed(03.1875,QstateIM(2)) then
				char2IM <= "+03.1875";
			elsif QstateIM(2) = to_sfixed(03.2500,QstateIM(2)) then
				char2IM <= "+03.2500";
			elsif QstateIM(2) = to_sfixed(03.3125,QstateIM(2)) then
				char2IM <= "+03.3125";
			elsif QstateIM(2) = to_sfixed(03.3750,QstateIM(2)) then
				char2IM <= "+03.3750";
			elsif QstateIM(2) = to_sfixed(03.4375,QstateIM(2)) then
				char2IM <= "+03.4375";
			elsif QstateIM(2) = to_sfixed(03.5000,QstateIM(2)) then
				char2IM <= "+03.5000";
			elsif QstateIM(2) = to_sfixed(03.5625,QstateIM(2)) then
				char2IM <= "+03.5625";
			elsif QstateIM(2) = to_sfixed(03.6250,QstateIM(2)) then
				char2IM <= "+03.6250";
			elsif QstateIM(2) = to_sfixed(03.6875,QstateIM(2)) then
				char2IM <= "+03.6875";
			elsif QstateIM(2) = to_sfixed(03.7500,QstateIM(2)) then
				char2IM <= "+03.7500";
			elsif QstateIM(2) = to_sfixed(03.8125,QstateIM(2)) then
				char2IM <= "+03.8125";
			elsif QstateIM(2) = to_sfixed(03.8750,QstateIM(2)) then
				char2IM <= "+03.8750";
			elsif QstateIM(2) = to_sfixed(03.9375,QstateIM(2)) then
				char2IM <= "+03.9375";
			elsif QstateIM(2) = to_sfixed(04.0000,QstateIM(2)) then
				char2IM <= "+04.0000";
			elsif QstateIM(2) = to_sfixed(04.0625,QstateIM(2)) then
				char2IM <= "+04.0625";
			elsif QstateIM(2) = to_sfixed(04.1250,QstateIM(2)) then
				char2IM <= "+04.1250";
			elsif QstateIM(2) = to_sfixed(04.1875,QstateIM(2)) then
				char2IM <= "+04.1875";
			elsif QstateIM(2) = to_sfixed(04.2500,QstateIM(2)) then
				char2IM <= "+04.2500";
			elsif QstateIM(2) = to_sfixed(04.3125,QstateIM(2)) then
				char2IM <= "+04.3125";
			elsif QstateIM(2) = to_sfixed(04.3750,QstateIM(2)) then
				char2IM <= "+04.3750";
			elsif QstateIM(2) = to_sfixed(04.4375,QstateIM(2)) then
				char2IM <= "+04.4375";
			elsif QstateIM(2) = to_sfixed(04.5000,QstateIM(2)) then
				char2IM <= "+04.5000";
			elsif QstateIM(2) = to_sfixed(04.5625,QstateIM(2)) then
				char2IM <= "+04.5625";
			elsif QstateIM(2) = to_sfixed(04.6250,QstateIM(2)) then
				char2IM <= "+04.6250";
			elsif QstateIM(2) = to_sfixed(04.6875,QstateIM(2)) then
				char2IM <= "+04.6875";
			elsif QstateIM(2) = to_sfixed(04.7500,QstateIM(2)) then
				char2IM <= "+04.7500";
			elsif QstateIM(2) = to_sfixed(04.8125,QstateIM(2)) then
				char2IM <= "+04.8125";
			elsif QstateIM(2) = to_sfixed(04.8750,QstateIM(2)) then
				char2IM <= "+04.8750";
			elsif QstateIM(2) = to_sfixed(04.9375,QstateIM(2)) then
				char2IM <= "+04.9375";
			elsif QstateIM(2) = to_sfixed(05.0000,QstateIM(2)) then
				char2IM <= "+05.0000";
			elsif QstateIM(2) = to_sfixed(05.0625,QstateIM(2)) then
				char2IM <= "+05.0625";
			elsif QstateIM(2) = to_sfixed(05.1250,QstateIM(2)) then
				char2IM <= "+05.1250";
			elsif QstateIM(2) = to_sfixed(05.1875,QstateIM(2)) then
				char2IM <= "+05.1875";
			elsif QstateIM(2) = to_sfixed(05.2500,QstateIM(2)) then
				char2IM <= "+05.2500";
			elsif QstateIM(2) = to_sfixed(05.3125,QstateIM(2)) then
				char2IM <= "+05.3125";
			elsif QstateIM(2) = to_sfixed(05.3750,QstateIM(2)) then
				char2IM <= "+05.3750";
			elsif QstateIM(2) = to_sfixed(05.4375,QstateIM(2)) then
				char2IM <= "+05.4375";
			elsif QstateIM(2) = to_sfixed(05.5000,QstateIM(2)) then
				char2IM <= "+05.5000";
			elsif QstateIM(2) = to_sfixed(05.5625,QstateIM(2)) then
				char2IM <= "+05.5625";
			elsif QstateIM(2) = to_sfixed(05.6250,QstateIM(2)) then
				char2IM <= "+05.6250";
			elsif QstateIM(2) = to_sfixed(05.6875,QstateIM(2)) then
				char2IM <= "+05.6875";
			elsif QstateIM(2) = to_sfixed(05.7500,QstateIM(2)) then
				char2IM <= "+05.7500";
			elsif QstateIM(2) = to_sfixed(05.8125,QstateIM(2)) then
				char2IM <= "+05.8125";
			elsif QstateIM(2) = to_sfixed(05.8750,QstateIM(2)) then
				char2IM <= "+05.8750";
			elsif QstateIM(2) = to_sfixed(05.9375,QstateIM(2)) then
				char2IM <= "+05.9375";
			elsif QstateIM(2) = to_sfixed(06.0000,QstateIM(2)) then
				char2IM <= "+06.0000";
			elsif QstateIM(2) = to_sfixed(06.0625,QstateIM(2)) then
				char2IM <= "+06.0625";
			elsif QstateIM(2) = to_sfixed(06.1250,QstateIM(2)) then
				char2IM <= "+06.1250";
			elsif QstateIM(2) = to_sfixed(06.1875,QstateIM(2)) then
				char2IM <= "+06.1875";
			elsif QstateIM(2) = to_sfixed(06.2500,QstateIM(2)) then
				char2IM <= "+06.2500";
			elsif QstateIM(2) = to_sfixed(06.3125,QstateIM(2)) then
				char2IM <= "+06.3125";
			elsif QstateIM(2) = to_sfixed(06.3750,QstateIM(2)) then
				char2IM <= "+06.3750";
			elsif QstateIM(2) = to_sfixed(06.4375,QstateIM(2)) then
				char2IM <= "+06.4375";
			elsif QstateIM(2) = to_sfixed(06.5000,QstateIM(2)) then
				char2IM <= "+06.5000";
			elsif QstateIM(2) = to_sfixed(06.5625,QstateIM(2)) then
				char2IM <= "+06.5625";
			elsif QstateIM(2) = to_sfixed(06.6250,QstateIM(2)) then
				char2IM <= "+06.6250";
			elsif QstateIM(2) = to_sfixed(06.6875,QstateIM(2)) then
				char2IM <= "+06.6875";
			elsif QstateIM(2) = to_sfixed(06.7500,QstateIM(2)) then
				char2IM <= "+06.7500";
			elsif QstateIM(2) = to_sfixed(06.8125,QstateIM(2)) then
				char2IM <= "+06.8125";
			elsif QstateIM(2) = to_sfixed(06.8750,QstateIM(2)) then
				char2IM <= "+06.8750";
			elsif QstateIM(2) = to_sfixed(06.9375,QstateIM(2)) then
				char2IM <= "+06.9375";
			elsif QstateIM(2) = to_sfixed(07.0000,QstateIM(2)) then
				char2IM <= "+07.0000";
			elsif QstateIM(2) = to_sfixed(07.0625,QstateIM(2)) then
				char2IM <= "+07.0625";
			elsif QstateIM(2) = to_sfixed(07.1250,QstateIM(2)) then
				char2IM <= "+07.1250";
			elsif QstateIM(2) = to_sfixed(07.1875,QstateIM(2)) then
				char2IM <= "+07.1875";
			elsif QstateIM(2) = to_sfixed(07.2500,QstateIM(2)) then
				char2IM <= "+07.2500";
			elsif QstateIM(2) = to_sfixed(07.3125,QstateIM(2)) then
				char2IM <= "+07.3125";
			elsif QstateIM(2) = to_sfixed(07.3750,QstateIM(2)) then
				char2IM <= "+07.3750";
			elsif QstateIM(2) = to_sfixed(07.4375,QstateIM(2)) then
				char2IM <= "+07.4375";
			elsif QstateIM(2) = to_sfixed(07.5000,QstateIM(2)) then
				char2IM <= "+07.5000";
			elsif QstateIM(2) = to_sfixed(07.5625,QstateIM(2)) then
				char2IM <= "+07.5625";
			elsif QstateIM(2) = to_sfixed(07.6250,QstateIM(2)) then
				char2IM <= "+07.6250";
			elsif QstateIM(2) = to_sfixed(07.6875,QstateIM(2)) then
				char2IM <= "+07.6875";
			elsif QstateIM(2) = to_sfixed(07.7500,QstateIM(2)) then
				char2IM <= "+07.7500";
			elsif QstateIM(2) = to_sfixed(07.8125,QstateIM(2)) then
				char2IM <= "+07.8125";
			elsif QstateIM(2) = to_sfixed(07.8750,QstateIM(2)) then
				char2IM <= "+07.8750";
			elsif QstateIM(2) = to_sfixed(07.9375,QstateIM(2)) then
				char2IM <= "+07.9375";
			elsif QstateIM(2) = to_sfixed(08.0000,QstateIM(2)) then
				char2IM <= "+08.0000";
			elsif QstateIM(2) = to_sfixed(08.0625,QstateIM(2)) then
				char2IM <= "+08.0625";
			elsif QstateIM(2) = to_sfixed(08.1250,QstateIM(2)) then
				char2IM <= "+08.1250";
			elsif QstateIM(2) = to_sfixed(08.1875,QstateIM(2)) then
				char2IM <= "+08.1875";
			elsif QstateIM(2) = to_sfixed(08.2500,QstateIM(2)) then
				char2IM <= "+08.2500";
			elsif QstateIM(2) = to_sfixed(08.3125,QstateIM(2)) then
				char2IM <= "+08.3125";
			elsif QstateIM(2) = to_sfixed(08.3750,QstateIM(2)) then
				char2IM <= "+08.3750";
			elsif QstateIM(2) = to_sfixed(08.4375,QstateIM(2)) then
				char2IM <= "+08.4375";
			elsif QstateIM(2) = to_sfixed(08.5000,QstateIM(2)) then
				char2IM <= "+08.5000";
			elsif QstateIM(2) = to_sfixed(08.5625,QstateIM(2)) then
				char2IM <= "+08.5625";
			elsif QstateIM(2) = to_sfixed(08.6250,QstateIM(2)) then
				char2IM <= "+08.6250";
			elsif QstateIM(2) = to_sfixed(08.6875,QstateIM(2)) then
				char2IM <= "+08.6875";
			elsif QstateIM(2) = to_sfixed(08.7500,QstateIM(2)) then
				char2IM <= "+08.7500";
			elsif QstateIM(2) = to_sfixed(08.8125,QstateIM(2)) then
				char2IM <= "+08.8125";
			elsif QstateIM(2) = to_sfixed(08.8750,QstateIM(2)) then
				char2IM <= "+08.8750";
			elsif QstateIM(2) = to_sfixed(08.9375,QstateIM(2)) then
				char2IM <= "+08.9375";
			elsif QstateIM(2) = to_sfixed(09.0000,QstateIM(2)) then
				char2IM <= "+09.0000";
			elsif QstateIM(2) = to_sfixed(09.0625,QstateIM(2)) then
				char2IM <= "+09.0625";
			elsif QstateIM(2) = to_sfixed(09.1250,QstateIM(2)) then
				char2IM <= "+09.1250";
			elsif QstateIM(2) = to_sfixed(09.1875,QstateIM(2)) then
				char2IM <= "+09.1875";
			elsif QstateIM(2) = to_sfixed(09.2500,QstateIM(2)) then
				char2IM <= "+09.2500";
			elsif QstateIM(2) = to_sfixed(09.3125,QstateIM(2)) then
				char2IM <= "+09.3125";
			elsif QstateIM(2) = to_sfixed(09.3750,QstateIM(2)) then
				char2IM <= "+09.3750";
			elsif QstateIM(2) = to_sfixed(09.4375,QstateIM(2)) then
				char2IM <= "+09.4375";
			elsif QstateIM(2) = to_sfixed(09.5000,QstateIM(2)) then
				char2IM <= "+09.5000";
			elsif QstateIM(2) = to_sfixed(09.5625,QstateIM(2)) then
				char2IM <= "+09.5625";
			elsif QstateIM(2) = to_sfixed(09.6250,QstateIM(2)) then
				char2IM <= "+09.6250";
			elsif QstateIM(2) = to_sfixed(09.6875,QstateIM(2)) then
				char2IM <= "+09.6875";
			elsif QstateIM(2) = to_sfixed(09.7500,QstateIM(2)) then
				char2IM <= "+09.7500";
			elsif QstateIM(2) = to_sfixed(09.8125,QstateIM(2)) then
				char2IM <= "+09.8125";
			elsif QstateIM(2) = to_sfixed(09.8750,QstateIM(2)) then
				char2IM <= "+09.8750";
			elsif QstateIM(2) = to_sfixed(09.9375,QstateIM(2)) then
				char2IM <= "+09.9375";
			elsif QstateIM(2) = to_sfixed(10.0000,QstateIM(2)) then
				char2IM <= "+10.0000";
			elsif QstateIM(2) = to_sfixed(10.0625,QstateIM(2)) then
				char2IM <= "+10.0625";
			elsif QstateIM(2) = to_sfixed(10.1250,QstateIM(2)) then
				char2IM <= "+10.1250";
			elsif QstateIM(2) = to_sfixed(10.1875,QstateIM(2)) then
				char2IM <= "+10.1875";
			elsif QstateIM(2) = to_sfixed(10.2500,QstateIM(2)) then
				char2IM <= "+10.2500";
			elsif QstateIM(2) = to_sfixed(10.3125,QstateIM(2)) then
				char2IM <= "+10.3125";
			elsif QstateIM(2) = to_sfixed(10.3750,QstateIM(2)) then
				char2IM <= "+10.3750";
			elsif QstateIM(2) = to_sfixed(10.4375,QstateIM(2)) then
				char2IM <= "+10.4375";
			elsif QstateIM(2) = to_sfixed(10.5000,QstateIM(2)) then
				char2IM <= "+10.5000";
			elsif QstateIM(2) = to_sfixed(10.5625,QstateIM(2)) then
				char2IM <= "+10.5625";
			elsif QstateIM(2) = to_sfixed(10.6250,QstateIM(2)) then
				char2IM <= "+10.6250";
			elsif QstateIM(2) = to_sfixed(10.6875,QstateIM(2)) then
				char2IM <= "+10.6875";
			elsif QstateIM(2) = to_sfixed(10.7500,QstateIM(2)) then
				char2IM <= "+10.7500";
			elsif QstateIM(2) = to_sfixed(10.8125,QstateIM(2)) then
				char2IM <= "+10.8125";
			elsif QstateIM(2) = to_sfixed(10.8750,QstateIM(2)) then
				char2IM <= "+10.8750";
			elsif QstateIM(2) = to_sfixed(10.9375,QstateIM(2)) then
				char2IM <= "+10.9375";
			elsif QstateIM(2) = to_sfixed(11.0000,QstateIM(2)) then
				char2IM <= "+11.0000";
			elsif QstateIM(2) = to_sfixed(11.0625,QstateIM(2)) then
				char2IM <= "+11.0625";
			elsif QstateIM(2) = to_sfixed(11.1250,QstateIM(2)) then
				char2IM <= "+11.1250";
			elsif QstateIM(2) = to_sfixed(11.1875,QstateIM(2)) then
				char2IM <= "+11.1875";
			elsif QstateIM(2) = to_sfixed(11.2500,QstateIM(2)) then
				char2IM <= "+11.2500";
			elsif QstateIM(2) = to_sfixed(11.3125,QstateIM(2)) then
				char2IM <= "+11.3125";
			elsif QstateIM(2) = to_sfixed(11.3750,QstateIM(2)) then
				char2IM <= "+11.3750";
			elsif QstateIM(2) = to_sfixed(11.4375,QstateIM(2)) then
				char2IM <= "+11.4375";
			elsif QstateIM(2) = to_sfixed(11.5000,QstateIM(2)) then
				char2IM <= "+11.5000";
			elsif QstateIM(2) = to_sfixed(11.5625,QstateIM(2)) then
				char2IM <= "+11.5625";
			elsif QstateIM(2) = to_sfixed(11.6250,QstateIM(2)) then
				char2IM <= "+11.6250";
			elsif QstateIM(2) = to_sfixed(11.6875,QstateIM(2)) then
				char2IM <= "+11.6875";
			elsif QstateIM(2) = to_sfixed(11.7500,QstateIM(2)) then
				char2IM <= "+11.7500";
			elsif QstateIM(2) = to_sfixed(11.8125,QstateIM(2)) then
				char2IM <= "+11.8125";
			elsif QstateIM(2) = to_sfixed(11.8750,QstateIM(2)) then
				char2IM <= "+11.8750";
			elsif QstateIM(2) = to_sfixed(11.9375,QstateIM(2)) then
				char2IM <= "+11.9375";
			elsif QstateIM(2) = to_sfixed(12.0000,QstateIM(2)) then
				char2IM <= "+12.0000";
			elsif QstateIM(2) = to_sfixed(12.0625,QstateIM(2)) then
				char2IM <= "+12.0625";
			elsif QstateIM(2) = to_sfixed(12.1250,QstateIM(2)) then
				char2IM <= "+12.1250";
			elsif QstateIM(2) = to_sfixed(12.1875,QstateIM(2)) then
				char2IM <= "+12.1875";
			elsif QstateIM(2) = to_sfixed(12.2500,QstateIM(2)) then
				char2IM <= "+12.2500";
			elsif QstateIM(2) = to_sfixed(12.3125,QstateIM(2)) then
				char2IM <= "+12.3125";
			elsif QstateIM(2) = to_sfixed(12.3750,QstateIM(2)) then
				char2IM <= "+12.3750";
			elsif QstateIM(2) = to_sfixed(12.4375,QstateIM(2)) then
				char2IM <= "+12.4375";
			elsif QstateIM(2) = to_sfixed(12.5000,QstateIM(2)) then
				char2IM <= "+12.5000";
			elsif QstateIM(2) = to_sfixed(12.5625,QstateIM(2)) then
				char2IM <= "+12.5625";
			elsif QstateIM(2) = to_sfixed(12.6250,QstateIM(2)) then
				char2IM <= "+12.6250";
			elsif QstateIM(2) = to_sfixed(12.6875,QstateIM(2)) then
				char2IM <= "+12.6875";
			elsif QstateIM(2) = to_sfixed(12.7500,QstateIM(2)) then
				char2IM <= "+12.7500";
			elsif QstateIM(2) = to_sfixed(12.8125,QstateIM(2)) then
				char2IM <= "+12.8125";
			elsif QstateIM(2) = to_sfixed(12.8750,QstateIM(2)) then
				char2IM <= "+12.8750";
			elsif QstateIM(2) = to_sfixed(12.9375,QstateIM(2)) then
				char2IM <= "+12.9375";
			elsif QstateIM(2) = to_sfixed(13.0000,QstateIM(2)) then
				char2IM <= "+13.0000";
			elsif QstateIM(2) = to_sfixed(13.0625,QstateIM(2)) then
				char2IM <= "+13.0625";
			elsif QstateIM(2) = to_sfixed(13.1250,QstateIM(2)) then
				char2IM <= "+13.1250";
			elsif QstateIM(2) = to_sfixed(13.1875,QstateIM(2)) then
				char2IM <= "+13.1875";
			elsif QstateIM(2) = to_sfixed(13.2500,QstateIM(2)) then
				char2IM <= "+13.2500";
			elsif QstateIM(2) = to_sfixed(13.3125,QstateIM(2)) then
				char2IM <= "+13.3125";
			elsif QstateIM(2) = to_sfixed(13.3750,QstateIM(2)) then
				char2IM <= "+13.3750";
			elsif QstateIM(2) = to_sfixed(13.4375,QstateIM(2)) then
				char2IM <= "+13.4375";
			elsif QstateIM(2) = to_sfixed(13.5000,QstateIM(2)) then
				char2IM <= "+13.5000";
			elsif QstateIM(2) = to_sfixed(13.5625,QstateIM(2)) then
				char2IM <= "+13.5625";
			elsif QstateIM(2) = to_sfixed(13.6250,QstateIM(2)) then
				char2IM <= "+13.6250";
			elsif QstateIM(2) = to_sfixed(13.6875,QstateIM(2)) then
				char2IM <= "+13.6875";
			elsif QstateIM(2) = to_sfixed(13.7500,QstateIM(2)) then
				char2IM <= "+13.7500";
			elsif QstateIM(2) = to_sfixed(13.8125,QstateIM(2)) then
				char2IM <= "+13.8125";
			elsif QstateIM(2) = to_sfixed(13.8750,QstateIM(2)) then
				char2IM <= "+13.8750";
			elsif QstateIM(2) = to_sfixed(13.9375,QstateIM(2)) then
				char2IM <= "+13.9375";
			elsif QstateIM(2) = to_sfixed(14.0000,QstateIM(2)) then
				char2IM <= "+14.0000";
			elsif QstateIM(2) = to_sfixed(14.0625,QstateIM(2)) then
				char2IM <= "+14.0625";
			elsif QstateIM(2) = to_sfixed(14.1250,QstateIM(2)) then
				char2IM <= "+14.1250";
			elsif QstateIM(2) = to_sfixed(14.1875,QstateIM(2)) then
				char2IM <= "+14.1875";
			elsif QstateIM(2) = to_sfixed(14.2500,QstateIM(2)) then
				char2IM <= "+14.2500";
			elsif QstateIM(2) = to_sfixed(14.3125,QstateIM(2)) then
				char2IM <= "+14.3125";
			elsif QstateIM(2) = to_sfixed(14.3750,QstateIM(2)) then
				char2IM <= "+14.3750";
			elsif QstateIM(2) = to_sfixed(14.4375,QstateIM(2)) then
				char2IM <= "+14.4375";
			elsif QstateIM(2) = to_sfixed(14.5000,QstateIM(2)) then
				char2IM <= "+14.5000";
			elsif QstateIM(2) = to_sfixed(14.5625,QstateIM(2)) then
				char2IM <= "+14.5625";
			elsif QstateIM(2) = to_sfixed(14.6250,QstateIM(2)) then
				char2IM <= "+14.6250";
			elsif QstateIM(2) = to_sfixed(14.6875,QstateIM(2)) then
				char2IM <= "+14.6875";
			elsif QstateIM(2) = to_sfixed(14.7500,QstateIM(2)) then
				char2IM <= "+14.7500";
			elsif QstateIM(2) = to_sfixed(14.8125,QstateIM(2)) then
				char2IM <= "+14.8125";
			elsif QstateIM(2) = to_sfixed(14.8750,QstateIM(2)) then
				char2IM <= "+14.8750";
			elsif QstateIM(2) = to_sfixed(14.9375,QstateIM(2)) then
				char2IM <= "+14.9375";
			elsif QstateIM(2) = to_sfixed(15.0000,QstateIM(2)) then
				char2IM <= "+15.0000";
			elsif QstateIM(2) = to_sfixed(15.0625,QstateIM(2)) then
				char2IM <= "+15.0625";
			elsif QstateIM(2) = to_sfixed(15.1250,QstateIM(2)) then
				char2IM <= "+15.1250";
			elsif QstateIM(2) = to_sfixed(15.1875,QstateIM(2)) then
				char2IM <= "+15.1875";
			elsif QstateIM(2) = to_sfixed(15.2500,QstateIM(2)) then
				char2IM <= "+15.2500";
			elsif QstateIM(2) = to_sfixed(15.3125,QstateIM(2)) then
				char2IM <= "+15.3125";
			elsif QstateIM(2) = to_sfixed(15.3750,QstateIM(2)) then
				char2IM <= "+15.3750";
			elsif QstateIM(2) = to_sfixed(15.4375,QstateIM(2)) then
				char2IM <= "+15.4375";
			elsif QstateIM(2) = to_sfixed(15.5000,QstateIM(2)) then
				char2IM <= "+15.5000";
			elsif QstateIM(2) = to_sfixed(15.5625,QstateIM(2)) then
				char2IM <= "+15.5625";
			elsif QstateIM(2) = to_sfixed(15.6250,QstateIM(2)) then
				char2IM <= "+15.6250";
			elsif QstateIM(2) = to_sfixed(15.6875,QstateIM(2)) then
				char2IM <= "+15.6875";
			elsif QstateIM(2) = to_sfixed(15.7500,QstateIM(2)) then
				char2IM <= "+15.7500";
			elsif QstateIM(2) = to_sfixed(15.8125,QstateIM(2)) then
				char2IM <= "+15.8125";
			elsif QstateIM(2) = to_sfixed(15.8750,QstateIM(2)) then
				char2IM <= "+15.8750";
			elsif QstateIM(2) = to_sfixed(15.9375,QstateIM(2)) then
				char2IM <= "+15.9375";
			end if;
			if QstateRE(3) = to_sfixed(-15.9375,QstateRE(3)) then
				char3RE <= "-15.9375";
			elsif QstateRE(3) = to_sfixed(-15.8750,QstateRE(3)) then
				char3RE <= "-15.8750";
			elsif QstateRE(3) = to_sfixed(-15.8125,QstateRE(3)) then
				char3RE <= "-15.8125";
			elsif QstateRE(3) = to_sfixed(-15.7500,QstateRE(3)) then
				char3RE <= "-15.7500";
			elsif QstateRE(3) = to_sfixed(-15.6875,QstateRE(3)) then
				char3RE <= "-15.6875";
			elsif QstateRE(3) = to_sfixed(-15.6250,QstateRE(3)) then
				char3RE <= "-15.6250";
			elsif QstateRE(3) = to_sfixed(-15.5625,QstateRE(3)) then
				char3RE <= "-15.5625";
			elsif QstateRE(3) = to_sfixed(-15.5000,QstateRE(3)) then
				char3RE <= "-15.5000";
			elsif QstateRE(3) = to_sfixed(-15.4375,QstateRE(3)) then
				char3RE <= "-15.4375";
			elsif QstateRE(3) = to_sfixed(-15.3750,QstateRE(3)) then
				char3RE <= "-15.3750";
			elsif QstateRE(3) = to_sfixed(-15.3125,QstateRE(3)) then
				char3RE <= "-15.3125";
			elsif QstateRE(3) = to_sfixed(-15.2500,QstateRE(3)) then
				char3RE <= "-15.2500";
			elsif QstateRE(3) = to_sfixed(-15.1875,QstateRE(3)) then
				char3RE <= "-15.1875";
			elsif QstateRE(3) = to_sfixed(-15.1250,QstateRE(3)) then
				char3RE <= "-15.1250";
			elsif QstateRE(3) = to_sfixed(-15.0625,QstateRE(3)) then
				char3RE <= "-15.0625";
			elsif QstateRE(3) = to_sfixed(-15.0000,QstateRE(3)) then
				char3RE <= "-15.0000";
			elsif QstateRE(3) = to_sfixed(-14.9375,QstateRE(3)) then
				char3RE <= "-14.9375";
			elsif QstateRE(3) = to_sfixed(-14.8750,QstateRE(3)) then
				char3RE <= "-14.8750";
			elsif QstateRE(3) = to_sfixed(-14.8125,QstateRE(3)) then
				char3RE <= "-14.8125";
			elsif QstateRE(3) = to_sfixed(-14.7500,QstateRE(3)) then
				char3RE <= "-14.7500";
			elsif QstateRE(3) = to_sfixed(-14.6875,QstateRE(3)) then
				char3RE <= "-14.6875";
			elsif QstateRE(3) = to_sfixed(-14.6250,QstateRE(3)) then
				char3RE <= "-14.6250";
			elsif QstateRE(3) = to_sfixed(-14.5625,QstateRE(3)) then
				char3RE <= "-14.5625";
			elsif QstateRE(3) = to_sfixed(-14.5000,QstateRE(3)) then
				char3RE <= "-14.5000";
			elsif QstateRE(3) = to_sfixed(-14.4375,QstateRE(3)) then
				char3RE <= "-14.4375";
			elsif QstateRE(3) = to_sfixed(-14.3750,QstateRE(3)) then
				char3RE <= "-14.3750";
			elsif QstateRE(3) = to_sfixed(-14.3125,QstateRE(3)) then
				char3RE <= "-14.3125";
			elsif QstateRE(3) = to_sfixed(-14.2500,QstateRE(3)) then
				char3RE <= "-14.2500";
			elsif QstateRE(3) = to_sfixed(-14.1875,QstateRE(3)) then
				char3RE <= "-14.1875";
			elsif QstateRE(3) = to_sfixed(-14.1250,QstateRE(3)) then
				char3RE <= "-14.1250";
			elsif QstateRE(3) = to_sfixed(-14.0625,QstateRE(3)) then
				char3RE <= "-14.0625";
			elsif QstateRE(3) = to_sfixed(-14.0000,QstateRE(3)) then
				char3RE <= "-14.0000";
			elsif QstateRE(3) = to_sfixed(-13.9375,QstateRE(3)) then
				char3RE <= "-13.9375";
			elsif QstateRE(3) = to_sfixed(-13.8750,QstateRE(3)) then
				char3RE <= "-13.8750";
			elsif QstateRE(3) = to_sfixed(-13.8125,QstateRE(3)) then
				char3RE <= "-13.8125";
			elsif QstateRE(3) = to_sfixed(-13.7500,QstateRE(3)) then
				char3RE <= "-13.7500";
			elsif QstateRE(3) = to_sfixed(-13.6875,QstateRE(3)) then
				char3RE <= "-13.6875";
			elsif QstateRE(3) = to_sfixed(-13.6250,QstateRE(3)) then
				char3RE <= "-13.6250";
			elsif QstateRE(3) = to_sfixed(-13.5625,QstateRE(3)) then
				char3RE <= "-13.5625";
			elsif QstateRE(3) = to_sfixed(-13.5000,QstateRE(3)) then
				char3RE <= "-13.5000";
			elsif QstateRE(3) = to_sfixed(-13.4375,QstateRE(3)) then
				char3RE <= "-13.4375";
			elsif QstateRE(3) = to_sfixed(-13.3750,QstateRE(3)) then
				char3RE <= "-13.3750";
			elsif QstateRE(3) = to_sfixed(-13.3125,QstateRE(3)) then
				char3RE <= "-13.3125";
			elsif QstateRE(3) = to_sfixed(-13.2500,QstateRE(3)) then
				char3RE <= "-13.2500";
			elsif QstateRE(3) = to_sfixed(-13.1875,QstateRE(3)) then
				char3RE <= "-13.1875";
			elsif QstateRE(3) = to_sfixed(-13.1250,QstateRE(3)) then
				char3RE <= "-13.1250";
			elsif QstateRE(3) = to_sfixed(-13.0625,QstateRE(3)) then
				char3RE <= "-13.0625";
			elsif QstateRE(3) = to_sfixed(-13.0000,QstateRE(3)) then
				char3RE <= "-13.0000";
			elsif QstateRE(3) = to_sfixed(-12.9375,QstateRE(3)) then
				char3RE <= "-12.9375";
			elsif QstateRE(3) = to_sfixed(-12.8750,QstateRE(3)) then
				char3RE <= "-12.8750";
			elsif QstateRE(3) = to_sfixed(-12.8125,QstateRE(3)) then
				char3RE <= "-12.8125";
			elsif QstateRE(3) = to_sfixed(-12.7500,QstateRE(3)) then
				char3RE <= "-12.7500";
			elsif QstateRE(3) = to_sfixed(-12.6875,QstateRE(3)) then
				char3RE <= "-12.6875";
			elsif QstateRE(3) = to_sfixed(-12.6250,QstateRE(3)) then
				char3RE <= "-12.6250";
			elsif QstateRE(3) = to_sfixed(-12.5625,QstateRE(3)) then
				char3RE <= "-12.5625";
			elsif QstateRE(3) = to_sfixed(-12.5000,QstateRE(3)) then
				char3RE <= "-12.5000";
			elsif QstateRE(3) = to_sfixed(-12.4375,QstateRE(3)) then
				char3RE <= "-12.4375";
			elsif QstateRE(3) = to_sfixed(-12.3750,QstateRE(3)) then
				char3RE <= "-12.3750";
			elsif QstateRE(3) = to_sfixed(-12.3125,QstateRE(3)) then
				char3RE <= "-12.3125";
			elsif QstateRE(3) = to_sfixed(-12.2500,QstateRE(3)) then
				char3RE <= "-12.2500";
			elsif QstateRE(3) = to_sfixed(-12.1875,QstateRE(3)) then
				char3RE <= "-12.1875";
			elsif QstateRE(3) = to_sfixed(-12.1250,QstateRE(3)) then
				char3RE <= "-12.1250";
			elsif QstateRE(3) = to_sfixed(-12.0625,QstateRE(3)) then
				char3RE <= "-12.0625";
			elsif QstateRE(3) = to_sfixed(-12.0000,QstateRE(3)) then
				char3RE <= "-12.0000";
			elsif QstateRE(3) = to_sfixed(-11.9375,QstateRE(3)) then
				char3RE <= "-11.9375";
			elsif QstateRE(3) = to_sfixed(-11.8750,QstateRE(3)) then
				char3RE <= "-11.8750";
			elsif QstateRE(3) = to_sfixed(-11.8125,QstateRE(3)) then
				char3RE <= "-11.8125";
			elsif QstateRE(3) = to_sfixed(-11.7500,QstateRE(3)) then
				char3RE <= "-11.7500";
			elsif QstateRE(3) = to_sfixed(-11.6875,QstateRE(3)) then
				char3RE <= "-11.6875";
			elsif QstateRE(3) = to_sfixed(-11.6250,QstateRE(3)) then
				char3RE <= "-11.6250";
			elsif QstateRE(3) = to_sfixed(-11.5625,QstateRE(3)) then
				char3RE <= "-11.5625";
			elsif QstateRE(3) = to_sfixed(-11.5000,QstateRE(3)) then
				char3RE <= "-11.5000";
			elsif QstateRE(3) = to_sfixed(-11.4375,QstateRE(3)) then
				char3RE <= "-11.4375";
			elsif QstateRE(3) = to_sfixed(-11.3750,QstateRE(3)) then
				char3RE <= "-11.3750";
			elsif QstateRE(3) = to_sfixed(-11.3125,QstateRE(3)) then
				char3RE <= "-11.3125";
			elsif QstateRE(3) = to_sfixed(-11.2500,QstateRE(3)) then
				char3RE <= "-11.2500";
			elsif QstateRE(3) = to_sfixed(-11.1875,QstateRE(3)) then
				char3RE <= "-11.1875";
			elsif QstateRE(3) = to_sfixed(-11.1250,QstateRE(3)) then
				char3RE <= "-11.1250";
			elsif QstateRE(3) = to_sfixed(-11.0625,QstateRE(3)) then
				char3RE <= "-11.0625";
			elsif QstateRE(3) = to_sfixed(-11.0000,QstateRE(3)) then
				char3RE <= "-11.0000";
			elsif QstateRE(3) = to_sfixed(-10.9375,QstateRE(3)) then
				char3RE <= "-10.9375";
			elsif QstateRE(3) = to_sfixed(-10.8750,QstateRE(3)) then
				char3RE <= "-10.8750";
			elsif QstateRE(3) = to_sfixed(-10.8125,QstateRE(3)) then
				char3RE <= "-10.8125";
			elsif QstateRE(3) = to_sfixed(-10.7500,QstateRE(3)) then
				char3RE <= "-10.7500";
			elsif QstateRE(3) = to_sfixed(-10.6875,QstateRE(3)) then
				char3RE <= "-10.6875";
			elsif QstateRE(3) = to_sfixed(-10.6250,QstateRE(3)) then
				char3RE <= "-10.6250";
			elsif QstateRE(3) = to_sfixed(-10.5625,QstateRE(3)) then
				char3RE <= "-10.5625";
			elsif QstateRE(3) = to_sfixed(-10.5000,QstateRE(3)) then
				char3RE <= "-10.5000";
			elsif QstateRE(3) = to_sfixed(-10.4375,QstateRE(3)) then
				char3RE <= "-10.4375";
			elsif QstateRE(3) = to_sfixed(-10.3750,QstateRE(3)) then
				char3RE <= "-10.3750";
			elsif QstateRE(3) = to_sfixed(-10.3125,QstateRE(3)) then
				char3RE <= "-10.3125";
			elsif QstateRE(3) = to_sfixed(-10.2500,QstateRE(3)) then
				char3RE <= "-10.2500";
			elsif QstateRE(3) = to_sfixed(-10.1875,QstateRE(3)) then
				char3RE <= "-10.1875";
			elsif QstateRE(3) = to_sfixed(-10.1250,QstateRE(3)) then
				char3RE <= "-10.1250";
			elsif QstateRE(3) = to_sfixed(-10.0625,QstateRE(3)) then
				char3RE <= "-10.0625";
			elsif QstateRE(3) = to_sfixed(-10.0000,QstateRE(3)) then
				char3RE <= "-10.0000";
			elsif QstateRE(3) = to_sfixed(-9.9375,QstateRE(3)) then
				char3RE <= "--9.9375";
			elsif QstateRE(3) = to_sfixed(-9.8750,QstateRE(3)) then
				char3RE <= "--9.8750";
			elsif QstateRE(3) = to_sfixed(-9.8125,QstateRE(3)) then
				char3RE <= "--9.8125";
			elsif QstateRE(3) = to_sfixed(-9.7500,QstateRE(3)) then
				char3RE <= "--9.7500";
			elsif QstateRE(3) = to_sfixed(-9.6875,QstateRE(3)) then
				char3RE <= "--9.6875";
			elsif QstateRE(3) = to_sfixed(-9.6250,QstateRE(3)) then
				char3RE <= "--9.6250";
			elsif QstateRE(3) = to_sfixed(-9.5625,QstateRE(3)) then
				char3RE <= "--9.5625";
			elsif QstateRE(3) = to_sfixed(-9.5000,QstateRE(3)) then
				char3RE <= "--9.5000";
			elsif QstateRE(3) = to_sfixed(-9.4375,QstateRE(3)) then
				char3RE <= "--9.4375";
			elsif QstateRE(3) = to_sfixed(-9.3750,QstateRE(3)) then
				char3RE <= "--9.3750";
			elsif QstateRE(3) = to_sfixed(-9.3125,QstateRE(3)) then
				char3RE <= "--9.3125";
			elsif QstateRE(3) = to_sfixed(-9.2500,QstateRE(3)) then
				char3RE <= "--9.2500";
			elsif QstateRE(3) = to_sfixed(-9.1875,QstateRE(3)) then
				char3RE <= "--9.1875";
			elsif QstateRE(3) = to_sfixed(-9.1250,QstateRE(3)) then
				char3RE <= "--9.1250";
			elsif QstateRE(3) = to_sfixed(-9.0625,QstateRE(3)) then
				char3RE <= "--9.0625";
			elsif QstateRE(3) = to_sfixed(-9.0000,QstateRE(3)) then
				char3RE <= "--9.0000";
			elsif QstateRE(3) = to_sfixed(-8.9375,QstateRE(3)) then
				char3RE <= "--8.9375";
			elsif QstateRE(3) = to_sfixed(-8.8750,QstateRE(3)) then
				char3RE <= "--8.8750";
			elsif QstateRE(3) = to_sfixed(-8.8125,QstateRE(3)) then
				char3RE <= "--8.8125";
			elsif QstateRE(3) = to_sfixed(-8.7500,QstateRE(3)) then
				char3RE <= "--8.7500";
			elsif QstateRE(3) = to_sfixed(-8.6875,QstateRE(3)) then
				char3RE <= "--8.6875";
			elsif QstateRE(3) = to_sfixed(-8.6250,QstateRE(3)) then
				char3RE <= "--8.6250";
			elsif QstateRE(3) = to_sfixed(-8.5625,QstateRE(3)) then
				char3RE <= "--8.5625";
			elsif QstateRE(3) = to_sfixed(-8.5000,QstateRE(3)) then
				char3RE <= "--8.5000";
			elsif QstateRE(3) = to_sfixed(-8.4375,QstateRE(3)) then
				char3RE <= "--8.4375";
			elsif QstateRE(3) = to_sfixed(-8.3750,QstateRE(3)) then
				char3RE <= "--8.3750";
			elsif QstateRE(3) = to_sfixed(-8.3125,QstateRE(3)) then
				char3RE <= "--8.3125";
			elsif QstateRE(3) = to_sfixed(-8.2500,QstateRE(3)) then
				char3RE <= "--8.2500";
			elsif QstateRE(3) = to_sfixed(-8.1875,QstateRE(3)) then
				char3RE <= "--8.1875";
			elsif QstateRE(3) = to_sfixed(-8.1250,QstateRE(3)) then
				char3RE <= "--8.1250";
			elsif QstateRE(3) = to_sfixed(-8.0625,QstateRE(3)) then
				char3RE <= "--8.0625";
			elsif QstateRE(3) = to_sfixed(-8.0000,QstateRE(3)) then
				char3RE <= "--8.0000";
			elsif QstateRE(3) = to_sfixed(-7.9375,QstateRE(3)) then
				char3RE <= "--7.9375";
			elsif QstateRE(3) = to_sfixed(-7.8750,QstateRE(3)) then
				char3RE <= "--7.8750";
			elsif QstateRE(3) = to_sfixed(-7.8125,QstateRE(3)) then
				char3RE <= "--7.8125";
			elsif QstateRE(3) = to_sfixed(-7.7500,QstateRE(3)) then
				char3RE <= "--7.7500";
			elsif QstateRE(3) = to_sfixed(-7.6875,QstateRE(3)) then
				char3RE <= "--7.6875";
			elsif QstateRE(3) = to_sfixed(-7.6250,QstateRE(3)) then
				char3RE <= "--7.6250";
			elsif QstateRE(3) = to_sfixed(-7.5625,QstateRE(3)) then
				char3RE <= "--7.5625";
			elsif QstateRE(3) = to_sfixed(-7.5000,QstateRE(3)) then
				char3RE <= "--7.5000";
			elsif QstateRE(3) = to_sfixed(-7.4375,QstateRE(3)) then
				char3RE <= "--7.4375";
			elsif QstateRE(3) = to_sfixed(-7.3750,QstateRE(3)) then
				char3RE <= "--7.3750";
			elsif QstateRE(3) = to_sfixed(-7.3125,QstateRE(3)) then
				char3RE <= "--7.3125";
			elsif QstateRE(3) = to_sfixed(-7.2500,QstateRE(3)) then
				char3RE <= "--7.2500";
			elsif QstateRE(3) = to_sfixed(-7.1875,QstateRE(3)) then
				char3RE <= "--7.1875";
			elsif QstateRE(3) = to_sfixed(-7.1250,QstateRE(3)) then
				char3RE <= "--7.1250";
			elsif QstateRE(3) = to_sfixed(-7.0625,QstateRE(3)) then
				char3RE <= "--7.0625";
			elsif QstateRE(3) = to_sfixed(-7.0000,QstateRE(3)) then
				char3RE <= "--7.0000";
			elsif QstateRE(3) = to_sfixed(-6.9375,QstateRE(3)) then
				char3RE <= "--6.9375";
			elsif QstateRE(3) = to_sfixed(-6.8750,QstateRE(3)) then
				char3RE <= "--6.8750";
			elsif QstateRE(3) = to_sfixed(-6.8125,QstateRE(3)) then
				char3RE <= "--6.8125";
			elsif QstateRE(3) = to_sfixed(-6.7500,QstateRE(3)) then
				char3RE <= "--6.7500";
			elsif QstateRE(3) = to_sfixed(-6.6875,QstateRE(3)) then
				char3RE <= "--6.6875";
			elsif QstateRE(3) = to_sfixed(-6.6250,QstateRE(3)) then
				char3RE <= "--6.6250";
			elsif QstateRE(3) = to_sfixed(-6.5625,QstateRE(3)) then
				char3RE <= "--6.5625";
			elsif QstateRE(3) = to_sfixed(-6.5000,QstateRE(3)) then
				char3RE <= "--6.5000";
			elsif QstateRE(3) = to_sfixed(-6.4375,QstateRE(3)) then
				char3RE <= "--6.4375";
			elsif QstateRE(3) = to_sfixed(-6.3750,QstateRE(3)) then
				char3RE <= "--6.3750";
			elsif QstateRE(3) = to_sfixed(-6.3125,QstateRE(3)) then
				char3RE <= "--6.3125";
			elsif QstateRE(3) = to_sfixed(-6.2500,QstateRE(3)) then
				char3RE <= "--6.2500";
			elsif QstateRE(3) = to_sfixed(-6.1875,QstateRE(3)) then
				char3RE <= "--6.1875";
			elsif QstateRE(3) = to_sfixed(-6.1250,QstateRE(3)) then
				char3RE <= "--6.1250";
			elsif QstateRE(3) = to_sfixed(-6.0625,QstateRE(3)) then
				char3RE <= "--6.0625";
			elsif QstateRE(3) = to_sfixed(-6.0000,QstateRE(3)) then
				char3RE <= "--6.0000";
			elsif QstateRE(3) = to_sfixed(-5.9375,QstateRE(3)) then
				char3RE <= "--5.9375";
			elsif QstateRE(3) = to_sfixed(-5.8750,QstateRE(3)) then
				char3RE <= "--5.8750";
			elsif QstateRE(3) = to_sfixed(-5.8125,QstateRE(3)) then
				char3RE <= "--5.8125";
			elsif QstateRE(3) = to_sfixed(-5.7500,QstateRE(3)) then
				char3RE <= "--5.7500";
			elsif QstateRE(3) = to_sfixed(-5.6875,QstateRE(3)) then
				char3RE <= "--5.6875";
			elsif QstateRE(3) = to_sfixed(-5.6250,QstateRE(3)) then
				char3RE <= "--5.6250";
			elsif QstateRE(3) = to_sfixed(-5.5625,QstateRE(3)) then
				char3RE <= "--5.5625";
			elsif QstateRE(3) = to_sfixed(-5.5000,QstateRE(3)) then
				char3RE <= "--5.5000";
			elsif QstateRE(3) = to_sfixed(-5.4375,QstateRE(3)) then
				char3RE <= "--5.4375";
			elsif QstateRE(3) = to_sfixed(-5.3750,QstateRE(3)) then
				char3RE <= "--5.3750";
			elsif QstateRE(3) = to_sfixed(-5.3125,QstateRE(3)) then
				char3RE <= "--5.3125";
			elsif QstateRE(3) = to_sfixed(-5.2500,QstateRE(3)) then
				char3RE <= "--5.2500";
			elsif QstateRE(3) = to_sfixed(-5.1875,QstateRE(3)) then
				char3RE <= "--5.1875";
			elsif QstateRE(3) = to_sfixed(-5.1250,QstateRE(3)) then
				char3RE <= "--5.1250";
			elsif QstateRE(3) = to_sfixed(-5.0625,QstateRE(3)) then
				char3RE <= "--5.0625";
			elsif QstateRE(3) = to_sfixed(-5.0000,QstateRE(3)) then
				char3RE <= "--5.0000";
			elsif QstateRE(3) = to_sfixed(-4.9375,QstateRE(3)) then
				char3RE <= "--4.9375";
			elsif QstateRE(3) = to_sfixed(-4.8750,QstateRE(3)) then
				char3RE <= "--4.8750";
			elsif QstateRE(3) = to_sfixed(-4.8125,QstateRE(3)) then
				char3RE <= "--4.8125";
			elsif QstateRE(3) = to_sfixed(-4.7500,QstateRE(3)) then
				char3RE <= "--4.7500";
			elsif QstateRE(3) = to_sfixed(-4.6875,QstateRE(3)) then
				char3RE <= "--4.6875";
			elsif QstateRE(3) = to_sfixed(-4.6250,QstateRE(3)) then
				char3RE <= "--4.6250";
			elsif QstateRE(3) = to_sfixed(-4.5625,QstateRE(3)) then
				char3RE <= "--4.5625";
			elsif QstateRE(3) = to_sfixed(-4.5000,QstateRE(3)) then
				char3RE <= "--4.5000";
			elsif QstateRE(3) = to_sfixed(-4.4375,QstateRE(3)) then
				char3RE <= "--4.4375";
			elsif QstateRE(3) = to_sfixed(-4.3750,QstateRE(3)) then
				char3RE <= "--4.3750";
			elsif QstateRE(3) = to_sfixed(-4.3125,QstateRE(3)) then
				char3RE <= "--4.3125";
			elsif QstateRE(3) = to_sfixed(-4.2500,QstateRE(3)) then
				char3RE <= "--4.2500";
			elsif QstateRE(3) = to_sfixed(-4.1875,QstateRE(3)) then
				char3RE <= "--4.1875";
			elsif QstateRE(3) = to_sfixed(-4.1250,QstateRE(3)) then
				char3RE <= "--4.1250";
			elsif QstateRE(3) = to_sfixed(-4.0625,QstateRE(3)) then
				char3RE <= "--4.0625";
			elsif QstateRE(3) = to_sfixed(-4.0000,QstateRE(3)) then
				char3RE <= "--4.0000";
			elsif QstateRE(3) = to_sfixed(-3.9375,QstateRE(3)) then
				char3RE <= "--3.9375";
			elsif QstateRE(3) = to_sfixed(-3.8750,QstateRE(3)) then
				char3RE <= "--3.8750";
			elsif QstateRE(3) = to_sfixed(-3.8125,QstateRE(3)) then
				char3RE <= "--3.8125";
			elsif QstateRE(3) = to_sfixed(-3.7500,QstateRE(3)) then
				char3RE <= "--3.7500";
			elsif QstateRE(3) = to_sfixed(-3.6875,QstateRE(3)) then
				char3RE <= "--3.6875";
			elsif QstateRE(3) = to_sfixed(-3.6250,QstateRE(3)) then
				char3RE <= "--3.6250";
			elsif QstateRE(3) = to_sfixed(-3.5625,QstateRE(3)) then
				char3RE <= "--3.5625";
			elsif QstateRE(3) = to_sfixed(-3.5000,QstateRE(3)) then
				char3RE <= "--3.5000";
			elsif QstateRE(3) = to_sfixed(-3.4375,QstateRE(3)) then
				char3RE <= "--3.4375";
			elsif QstateRE(3) = to_sfixed(-3.3750,QstateRE(3)) then
				char3RE <= "--3.3750";
			elsif QstateRE(3) = to_sfixed(-3.3125,QstateRE(3)) then
				char3RE <= "--3.3125";
			elsif QstateRE(3) = to_sfixed(-3.2500,QstateRE(3)) then
				char3RE <= "--3.2500";
			elsif QstateRE(3) = to_sfixed(-3.1875,QstateRE(3)) then
				char3RE <= "--3.1875";
			elsif QstateRE(3) = to_sfixed(-3.1250,QstateRE(3)) then
				char3RE <= "--3.1250";
			elsif QstateRE(3) = to_sfixed(-3.0625,QstateRE(3)) then
				char3RE <= "--3.0625";
			elsif QstateRE(3) = to_sfixed(-3.0000,QstateRE(3)) then
				char3RE <= "--3.0000";
			elsif QstateRE(3) = to_sfixed(-2.9375,QstateRE(3)) then
				char3RE <= "--2.9375";
			elsif QstateRE(3) = to_sfixed(-2.8750,QstateRE(3)) then
				char3RE <= "--2.8750";
			elsif QstateRE(3) = to_sfixed(-2.8125,QstateRE(3)) then
				char3RE <= "--2.8125";
			elsif QstateRE(3) = to_sfixed(-2.7500,QstateRE(3)) then
				char3RE <= "--2.7500";
			elsif QstateRE(3) = to_sfixed(-2.6875,QstateRE(3)) then
				char3RE <= "--2.6875";
			elsif QstateRE(3) = to_sfixed(-2.6250,QstateRE(3)) then
				char3RE <= "--2.6250";
			elsif QstateRE(3) = to_sfixed(-2.5625,QstateRE(3)) then
				char3RE <= "--2.5625";
			elsif QstateRE(3) = to_sfixed(-2.5000,QstateRE(3)) then
				char3RE <= "--2.5000";
			elsif QstateRE(3) = to_sfixed(-2.4375,QstateRE(3)) then
				char3RE <= "--2.4375";
			elsif QstateRE(3) = to_sfixed(-2.3750,QstateRE(3)) then
				char3RE <= "--2.3750";
			elsif QstateRE(3) = to_sfixed(-2.3125,QstateRE(3)) then
				char3RE <= "--2.3125";
			elsif QstateRE(3) = to_sfixed(-2.2500,QstateRE(3)) then
				char3RE <= "--2.2500";
			elsif QstateRE(3) = to_sfixed(-2.1875,QstateRE(3)) then
				char3RE <= "--2.1875";
			elsif QstateRE(3) = to_sfixed(-2.1250,QstateRE(3)) then
				char3RE <= "--2.1250";
			elsif QstateRE(3) = to_sfixed(-2.0625,QstateRE(3)) then
				char3RE <= "--2.0625";
			elsif QstateRE(3) = to_sfixed(-2.0000,QstateRE(3)) then
				char3RE <= "--2.0000";
			elsif QstateRE(3) = to_sfixed(-1.9375,QstateRE(3)) then
				char3RE <= "--1.9375";
			elsif QstateRE(3) = to_sfixed(-1.8750,QstateRE(3)) then
				char3RE <= "--1.8750";
			elsif QstateRE(3) = to_sfixed(-1.8125,QstateRE(3)) then
				char3RE <= "--1.8125";
			elsif QstateRE(3) = to_sfixed(-1.7500,QstateRE(3)) then
				char3RE <= "--1.7500";
			elsif QstateRE(3) = to_sfixed(-1.6875,QstateRE(3)) then
				char3RE <= "--1.6875";
			elsif QstateRE(3) = to_sfixed(-1.6250,QstateRE(3)) then
				char3RE <= "--1.6250";
			elsif QstateRE(3) = to_sfixed(-1.5625,QstateRE(3)) then
				char3RE <= "--1.5625";
			elsif QstateRE(3) = to_sfixed(-1.5000,QstateRE(3)) then
				char3RE <= "--1.5000";
			elsif QstateRE(3) = to_sfixed(-1.4375,QstateRE(3)) then
				char3RE <= "--1.4375";
			elsif QstateRE(3) = to_sfixed(-1.3750,QstateRE(3)) then
				char3RE <= "--1.3750";
			elsif QstateRE(3) = to_sfixed(-1.3125,QstateRE(3)) then
				char3RE <= "--1.3125";
			elsif QstateRE(3) = to_sfixed(-1.2500,QstateRE(3)) then
				char3RE <= "--1.2500";
			elsif QstateRE(3) = to_sfixed(-1.1875,QstateRE(3)) then
				char3RE <= "--1.1875";
			elsif QstateRE(3) = to_sfixed(-1.1250,QstateRE(3)) then
				char3RE <= "--1.1250";
			elsif QstateRE(3) = to_sfixed(-1.0625,QstateRE(3)) then
				char3RE <= "--1.0625";
			elsif QstateRE(3) = to_sfixed(-1.0000,QstateRE(3)) then
				char3RE <= "--1.0000";
			elsif QstateRE(3) = to_sfixed(-0.9375,QstateRE(3)) then
				char3RE <= "--0.9375";
			elsif QstateRE(3) = to_sfixed(-0.8750,QstateRE(3)) then
				char3RE <= "--0.8750";
			elsif QstateRE(3) = to_sfixed(-0.8125,QstateRE(3)) then
				char3RE <= "--0.8125";
			elsif QstateRE(3) = to_sfixed(-0.7500,QstateRE(3)) then
				char3RE <= "--0.7500";
			elsif QstateRE(3) = to_sfixed(-0.6875,QstateRE(3)) then
				char3RE <= "--0.6875";
			elsif QstateRE(3) = to_sfixed(-0.6250,QstateRE(3)) then
				char3RE <= "--0.6250";
			elsif QstateRE(3) = to_sfixed(-0.5625,QstateRE(3)) then
				char3RE <= "--0.5625";
			elsif QstateRE(3) = to_sfixed(-0.5000,QstateRE(3)) then
				char3RE <= "--0.5000";
			elsif QstateRE(3) = to_sfixed(-0.4375,QstateRE(3)) then
				char3RE <= "--0.4375";
			elsif QstateRE(3) = to_sfixed(-0.3750,QstateRE(3)) then
				char3RE <= "--0.3750";
			elsif QstateRE(3) = to_sfixed(-0.3125,QstateRE(3)) then
				char3RE <= "--0.3125";
			elsif QstateRE(3) = to_sfixed(-0.2500,QstateRE(3)) then
				char3RE <= "--0.2500";
			elsif QstateRE(3) = to_sfixed(-0.1875,QstateRE(3)) then
				char3RE <= "--0.1875";
			elsif QstateRE(3) = to_sfixed(-0.1250,QstateRE(3)) then
				char3RE <= "--0.1250";
			elsif QstateRE(3) = to_sfixed(-0.0625,QstateRE(3)) then
				char3RE <= "--0.0625";
			elsif QstateRE(3) = to_sfixed(00.0000,QstateRE(3)) then
				char3RE <= "+00.0000";
			elsif QstateRE(3) = to_sfixed(00.0625,QstateRE(3)) then
				char3RE <= "+00.0625";
			elsif QstateRE(3) = to_sfixed(00.1250,QstateRE(3)) then
				char3RE <= "+00.1250";
			elsif QstateRE(3) = to_sfixed(00.1875,QstateRE(3)) then
				char3RE <= "+00.1875";
			elsif QstateRE(3) = to_sfixed(00.2500,QstateRE(3)) then
				char3RE <= "+00.2500";
			elsif QstateRE(3) = to_sfixed(00.3125,QstateRE(3)) then
				char3RE <= "+00.3125";
			elsif QstateRE(3) = to_sfixed(00.3750,QstateRE(3)) then
				char3RE <= "+00.3750";
			elsif QstateRE(3) = to_sfixed(00.4375,QstateRE(3)) then
				char3RE <= "+00.4375";
			elsif QstateRE(3) = to_sfixed(00.5000,QstateRE(3)) then
				char3RE <= "+00.5000";
			elsif QstateRE(3) = to_sfixed(00.5625,QstateRE(3)) then
				char3RE <= "+00.5625";
			elsif QstateRE(3) = to_sfixed(00.6250,QstateRE(3)) then
				char3RE <= "+00.6250";
			elsif QstateRE(3) = to_sfixed(00.6875,QstateRE(3)) then
				char3RE <= "+00.6875";
			elsif QstateRE(3) = to_sfixed(00.7500,QstateRE(3)) then
				char3RE <= "+00.7500";
			elsif QstateRE(3) = to_sfixed(00.8125,QstateRE(3)) then
				char3RE <= "+00.8125";
			elsif QstateRE(3) = to_sfixed(00.8750,QstateRE(3)) then
				char3RE <= "+00.8750";
			elsif QstateRE(3) = to_sfixed(00.9375,QstateRE(3)) then
				char3RE <= "+00.9375";
			elsif QstateRE(3) = to_sfixed(01.0000,QstateRE(3)) then
				char3RE <= "+01.0000";
			elsif QstateRE(3) = to_sfixed(01.0625,QstateRE(3)) then
				char3RE <= "+01.0625";
			elsif QstateRE(3) = to_sfixed(01.1250,QstateRE(3)) then
				char3RE <= "+01.1250";
			elsif QstateRE(3) = to_sfixed(01.1875,QstateRE(3)) then
				char3RE <= "+01.1875";
			elsif QstateRE(3) = to_sfixed(01.2500,QstateRE(3)) then
				char3RE <= "+01.2500";
			elsif QstateRE(3) = to_sfixed(01.3125,QstateRE(3)) then
				char3RE <= "+01.3125";
			elsif QstateRE(3) = to_sfixed(01.3750,QstateRE(3)) then
				char3RE <= "+01.3750";
			elsif QstateRE(3) = to_sfixed(01.4375,QstateRE(3)) then
				char3RE <= "+01.4375";
			elsif QstateRE(3) = to_sfixed(01.5000,QstateRE(3)) then
				char3RE <= "+01.5000";
			elsif QstateRE(3) = to_sfixed(01.5625,QstateRE(3)) then
				char3RE <= "+01.5625";
			elsif QstateRE(3) = to_sfixed(01.6250,QstateRE(3)) then
				char3RE <= "+01.6250";
			elsif QstateRE(3) = to_sfixed(01.6875,QstateRE(3)) then
				char3RE <= "+01.6875";
			elsif QstateRE(3) = to_sfixed(01.7500,QstateRE(3)) then
				char3RE <= "+01.7500";
			elsif QstateRE(3) = to_sfixed(01.8125,QstateRE(3)) then
				char3RE <= "+01.8125";
			elsif QstateRE(3) = to_sfixed(01.8750,QstateRE(3)) then
				char3RE <= "+01.8750";
			elsif QstateRE(3) = to_sfixed(01.9375,QstateRE(3)) then
				char3RE <= "+01.9375";
			elsif QstateRE(3) = to_sfixed(02.0000,QstateRE(3)) then
				char3RE <= "+02.0000";
			elsif QstateRE(3) = to_sfixed(02.0625,QstateRE(3)) then
				char3RE <= "+02.0625";
			elsif QstateRE(3) = to_sfixed(02.1250,QstateRE(3)) then
				char3RE <= "+02.1250";
			elsif QstateRE(3) = to_sfixed(02.1875,QstateRE(3)) then
				char3RE <= "+02.1875";
			elsif QstateRE(3) = to_sfixed(02.2500,QstateRE(3)) then
				char3RE <= "+02.2500";
			elsif QstateRE(3) = to_sfixed(02.3125,QstateRE(3)) then
				char3RE <= "+02.3125";
			elsif QstateRE(3) = to_sfixed(02.3750,QstateRE(3)) then
				char3RE <= "+02.3750";
			elsif QstateRE(3) = to_sfixed(02.4375,QstateRE(3)) then
				char3RE <= "+02.4375";
			elsif QstateRE(3) = to_sfixed(02.5000,QstateRE(3)) then
				char3RE <= "+02.5000";
			elsif QstateRE(3) = to_sfixed(02.5625,QstateRE(3)) then
				char3RE <= "+02.5625";
			elsif QstateRE(3) = to_sfixed(02.6250,QstateRE(3)) then
				char3RE <= "+02.6250";
			elsif QstateRE(3) = to_sfixed(02.6875,QstateRE(3)) then
				char3RE <= "+02.6875";
			elsif QstateRE(3) = to_sfixed(02.7500,QstateRE(3)) then
				char3RE <= "+02.7500";
			elsif QstateRE(3) = to_sfixed(02.8125,QstateRE(3)) then
				char3RE <= "+02.8125";
			elsif QstateRE(3) = to_sfixed(02.8750,QstateRE(3)) then
				char3RE <= "+02.8750";
			elsif QstateRE(3) = to_sfixed(02.9375,QstateRE(3)) then
				char3RE <= "+02.9375";
			elsif QstateRE(3) = to_sfixed(03.0000,QstateRE(3)) then
				char3RE <= "+03.0000";
			elsif QstateRE(3) = to_sfixed(03.0625,QstateRE(3)) then
				char3RE <= "+03.0625";
			elsif QstateRE(3) = to_sfixed(03.1250,QstateRE(3)) then
				char3RE <= "+03.1250";
			elsif QstateRE(3) = to_sfixed(03.1875,QstateRE(3)) then
				char3RE <= "+03.1875";
			elsif QstateRE(3) = to_sfixed(03.2500,QstateRE(3)) then
				char3RE <= "+03.2500";
			elsif QstateRE(3) = to_sfixed(03.3125,QstateRE(3)) then
				char3RE <= "+03.3125";
			elsif QstateRE(3) = to_sfixed(03.3750,QstateRE(3)) then
				char3RE <= "+03.3750";
			elsif QstateRE(3) = to_sfixed(03.4375,QstateRE(3)) then
				char3RE <= "+03.4375";
			elsif QstateRE(3) = to_sfixed(03.5000,QstateRE(3)) then
				char3RE <= "+03.5000";
			elsif QstateRE(3) = to_sfixed(03.5625,QstateRE(3)) then
				char3RE <= "+03.5625";
			elsif QstateRE(3) = to_sfixed(03.6250,QstateRE(3)) then
				char3RE <= "+03.6250";
			elsif QstateRE(3) = to_sfixed(03.6875,QstateRE(3)) then
				char3RE <= "+03.6875";
			elsif QstateRE(3) = to_sfixed(03.7500,QstateRE(3)) then
				char3RE <= "+03.7500";
			elsif QstateRE(3) = to_sfixed(03.8125,QstateRE(3)) then
				char3RE <= "+03.8125";
			elsif QstateRE(3) = to_sfixed(03.8750,QstateRE(3)) then
				char3RE <= "+03.8750";
			elsif QstateRE(3) = to_sfixed(03.9375,QstateRE(3)) then
				char3RE <= "+03.9375";
			elsif QstateRE(3) = to_sfixed(04.0000,QstateRE(3)) then
				char3RE <= "+04.0000";
			elsif QstateRE(3) = to_sfixed(04.0625,QstateRE(3)) then
				char3RE <= "+04.0625";
			elsif QstateRE(3) = to_sfixed(04.1250,QstateRE(3)) then
				char3RE <= "+04.1250";
			elsif QstateRE(3) = to_sfixed(04.1875,QstateRE(3)) then
				char3RE <= "+04.1875";
			elsif QstateRE(3) = to_sfixed(04.2500,QstateRE(3)) then
				char3RE <= "+04.2500";
			elsif QstateRE(3) = to_sfixed(04.3125,QstateRE(3)) then
				char3RE <= "+04.3125";
			elsif QstateRE(3) = to_sfixed(04.3750,QstateRE(3)) then
				char3RE <= "+04.3750";
			elsif QstateRE(3) = to_sfixed(04.4375,QstateRE(3)) then
				char3RE <= "+04.4375";
			elsif QstateRE(3) = to_sfixed(04.5000,QstateRE(3)) then
				char3RE <= "+04.5000";
			elsif QstateRE(3) = to_sfixed(04.5625,QstateRE(3)) then
				char3RE <= "+04.5625";
			elsif QstateRE(3) = to_sfixed(04.6250,QstateRE(3)) then
				char3RE <= "+04.6250";
			elsif QstateRE(3) = to_sfixed(04.6875,QstateRE(3)) then
				char3RE <= "+04.6875";
			elsif QstateRE(3) = to_sfixed(04.7500,QstateRE(3)) then
				char3RE <= "+04.7500";
			elsif QstateRE(3) = to_sfixed(04.8125,QstateRE(3)) then
				char3RE <= "+04.8125";
			elsif QstateRE(3) = to_sfixed(04.8750,QstateRE(3)) then
				char3RE <= "+04.8750";
			elsif QstateRE(3) = to_sfixed(04.9375,QstateRE(3)) then
				char3RE <= "+04.9375";
			elsif QstateRE(3) = to_sfixed(05.0000,QstateRE(3)) then
				char3RE <= "+05.0000";
			elsif QstateRE(3) = to_sfixed(05.0625,QstateRE(3)) then
				char3RE <= "+05.0625";
			elsif QstateRE(3) = to_sfixed(05.1250,QstateRE(3)) then
				char3RE <= "+05.1250";
			elsif QstateRE(3) = to_sfixed(05.1875,QstateRE(3)) then
				char3RE <= "+05.1875";
			elsif QstateRE(3) = to_sfixed(05.2500,QstateRE(3)) then
				char3RE <= "+05.2500";
			elsif QstateRE(3) = to_sfixed(05.3125,QstateRE(3)) then
				char3RE <= "+05.3125";
			elsif QstateRE(3) = to_sfixed(05.3750,QstateRE(3)) then
				char3RE <= "+05.3750";
			elsif QstateRE(3) = to_sfixed(05.4375,QstateRE(3)) then
				char3RE <= "+05.4375";
			elsif QstateRE(3) = to_sfixed(05.5000,QstateRE(3)) then
				char3RE <= "+05.5000";
			elsif QstateRE(3) = to_sfixed(05.5625,QstateRE(3)) then
				char3RE <= "+05.5625";
			elsif QstateRE(3) = to_sfixed(05.6250,QstateRE(3)) then
				char3RE <= "+05.6250";
			elsif QstateRE(3) = to_sfixed(05.6875,QstateRE(3)) then
				char3RE <= "+05.6875";
			elsif QstateRE(3) = to_sfixed(05.7500,QstateRE(3)) then
				char3RE <= "+05.7500";
			elsif QstateRE(3) = to_sfixed(05.8125,QstateRE(3)) then
				char3RE <= "+05.8125";
			elsif QstateRE(3) = to_sfixed(05.8750,QstateRE(3)) then
				char3RE <= "+05.8750";
			elsif QstateRE(3) = to_sfixed(05.9375,QstateRE(3)) then
				char3RE <= "+05.9375";
			elsif QstateRE(3) = to_sfixed(06.0000,QstateRE(3)) then
				char3RE <= "+06.0000";
			elsif QstateRE(3) = to_sfixed(06.0625,QstateRE(3)) then
				char3RE <= "+06.0625";
			elsif QstateRE(3) = to_sfixed(06.1250,QstateRE(3)) then
				char3RE <= "+06.1250";
			elsif QstateRE(3) = to_sfixed(06.1875,QstateRE(3)) then
				char3RE <= "+06.1875";
			elsif QstateRE(3) = to_sfixed(06.2500,QstateRE(3)) then
				char3RE <= "+06.2500";
			elsif QstateRE(3) = to_sfixed(06.3125,QstateRE(3)) then
				char3RE <= "+06.3125";
			elsif QstateRE(3) = to_sfixed(06.3750,QstateRE(3)) then
				char3RE <= "+06.3750";
			elsif QstateRE(3) = to_sfixed(06.4375,QstateRE(3)) then
				char3RE <= "+06.4375";
			elsif QstateRE(3) = to_sfixed(06.5000,QstateRE(3)) then
				char3RE <= "+06.5000";
			elsif QstateRE(3) = to_sfixed(06.5625,QstateRE(3)) then
				char3RE <= "+06.5625";
			elsif QstateRE(3) = to_sfixed(06.6250,QstateRE(3)) then
				char3RE <= "+06.6250";
			elsif QstateRE(3) = to_sfixed(06.6875,QstateRE(3)) then
				char3RE <= "+06.6875";
			elsif QstateRE(3) = to_sfixed(06.7500,QstateRE(3)) then
				char3RE <= "+06.7500";
			elsif QstateRE(3) = to_sfixed(06.8125,QstateRE(3)) then
				char3RE <= "+06.8125";
			elsif QstateRE(3) = to_sfixed(06.8750,QstateRE(3)) then
				char3RE <= "+06.8750";
			elsif QstateRE(3) = to_sfixed(06.9375,QstateRE(3)) then
				char3RE <= "+06.9375";
			elsif QstateRE(3) = to_sfixed(07.0000,QstateRE(3)) then
				char3RE <= "+07.0000";
			elsif QstateRE(3) = to_sfixed(07.0625,QstateRE(3)) then
				char3RE <= "+07.0625";
			elsif QstateRE(3) = to_sfixed(07.1250,QstateRE(3)) then
				char3RE <= "+07.1250";
			elsif QstateRE(3) = to_sfixed(07.1875,QstateRE(3)) then
				char3RE <= "+07.1875";
			elsif QstateRE(3) = to_sfixed(07.2500,QstateRE(3)) then
				char3RE <= "+07.2500";
			elsif QstateRE(3) = to_sfixed(07.3125,QstateRE(3)) then
				char3RE <= "+07.3125";
			elsif QstateRE(3) = to_sfixed(07.3750,QstateRE(3)) then
				char3RE <= "+07.3750";
			elsif QstateRE(3) = to_sfixed(07.4375,QstateRE(3)) then
				char3RE <= "+07.4375";
			elsif QstateRE(3) = to_sfixed(07.5000,QstateRE(3)) then
				char3RE <= "+07.5000";
			elsif QstateRE(3) = to_sfixed(07.5625,QstateRE(3)) then
				char3RE <= "+07.5625";
			elsif QstateRE(3) = to_sfixed(07.6250,QstateRE(3)) then
				char3RE <= "+07.6250";
			elsif QstateRE(3) = to_sfixed(07.6875,QstateRE(3)) then
				char3RE <= "+07.6875";
			elsif QstateRE(3) = to_sfixed(07.7500,QstateRE(3)) then
				char3RE <= "+07.7500";
			elsif QstateRE(3) = to_sfixed(07.8125,QstateRE(3)) then
				char3RE <= "+07.8125";
			elsif QstateRE(3) = to_sfixed(07.8750,QstateRE(3)) then
				char3RE <= "+07.8750";
			elsif QstateRE(3) = to_sfixed(07.9375,QstateRE(3)) then
				char3RE <= "+07.9375";
			elsif QstateRE(3) = to_sfixed(08.0000,QstateRE(3)) then
				char3RE <= "+08.0000";
			elsif QstateRE(3) = to_sfixed(08.0625,QstateRE(3)) then
				char3RE <= "+08.0625";
			elsif QstateRE(3) = to_sfixed(08.1250,QstateRE(3)) then
				char3RE <= "+08.1250";
			elsif QstateRE(3) = to_sfixed(08.1875,QstateRE(3)) then
				char3RE <= "+08.1875";
			elsif QstateRE(3) = to_sfixed(08.2500,QstateRE(3)) then
				char3RE <= "+08.2500";
			elsif QstateRE(3) = to_sfixed(08.3125,QstateRE(3)) then
				char3RE <= "+08.3125";
			elsif QstateRE(3) = to_sfixed(08.3750,QstateRE(3)) then
				char3RE <= "+08.3750";
			elsif QstateRE(3) = to_sfixed(08.4375,QstateRE(3)) then
				char3RE <= "+08.4375";
			elsif QstateRE(3) = to_sfixed(08.5000,QstateRE(3)) then
				char3RE <= "+08.5000";
			elsif QstateRE(3) = to_sfixed(08.5625,QstateRE(3)) then
				char3RE <= "+08.5625";
			elsif QstateRE(3) = to_sfixed(08.6250,QstateRE(3)) then
				char3RE <= "+08.6250";
			elsif QstateRE(3) = to_sfixed(08.6875,QstateRE(3)) then
				char3RE <= "+08.6875";
			elsif QstateRE(3) = to_sfixed(08.7500,QstateRE(3)) then
				char3RE <= "+08.7500";
			elsif QstateRE(3) = to_sfixed(08.8125,QstateRE(3)) then
				char3RE <= "+08.8125";
			elsif QstateRE(3) = to_sfixed(08.8750,QstateRE(3)) then
				char3RE <= "+08.8750";
			elsif QstateRE(3) = to_sfixed(08.9375,QstateRE(3)) then
				char3RE <= "+08.9375";
			elsif QstateRE(3) = to_sfixed(09.0000,QstateRE(3)) then
				char3RE <= "+09.0000";
			elsif QstateRE(3) = to_sfixed(09.0625,QstateRE(3)) then
				char3RE <= "+09.0625";
			elsif QstateRE(3) = to_sfixed(09.1250,QstateRE(3)) then
				char3RE <= "+09.1250";
			elsif QstateRE(3) = to_sfixed(09.1875,QstateRE(3)) then
				char3RE <= "+09.1875";
			elsif QstateRE(3) = to_sfixed(09.2500,QstateRE(3)) then
				char3RE <= "+09.2500";
			elsif QstateRE(3) = to_sfixed(09.3125,QstateRE(3)) then
				char3RE <= "+09.3125";
			elsif QstateRE(3) = to_sfixed(09.3750,QstateRE(3)) then
				char3RE <= "+09.3750";
			elsif QstateRE(3) = to_sfixed(09.4375,QstateRE(3)) then
				char3RE <= "+09.4375";
			elsif QstateRE(3) = to_sfixed(09.5000,QstateRE(3)) then
				char3RE <= "+09.5000";
			elsif QstateRE(3) = to_sfixed(09.5625,QstateRE(3)) then
				char3RE <= "+09.5625";
			elsif QstateRE(3) = to_sfixed(09.6250,QstateRE(3)) then
				char3RE <= "+09.6250";
			elsif QstateRE(3) = to_sfixed(09.6875,QstateRE(3)) then
				char3RE <= "+09.6875";
			elsif QstateRE(3) = to_sfixed(09.7500,QstateRE(3)) then
				char3RE <= "+09.7500";
			elsif QstateRE(3) = to_sfixed(09.8125,QstateRE(3)) then
				char3RE <= "+09.8125";
			elsif QstateRE(3) = to_sfixed(09.8750,QstateRE(3)) then
				char3RE <= "+09.8750";
			elsif QstateRE(3) = to_sfixed(09.9375,QstateRE(3)) then
				char3RE <= "+09.9375";
			elsif QstateRE(3) = to_sfixed(10.0000,QstateRE(3)) then
				char3RE <= "+10.0000";
			elsif QstateRE(3) = to_sfixed(10.0625,QstateRE(3)) then
				char3RE <= "+10.0625";
			elsif QstateRE(3) = to_sfixed(10.1250,QstateRE(3)) then
				char3RE <= "+10.1250";
			elsif QstateRE(3) = to_sfixed(10.1875,QstateRE(3)) then
				char3RE <= "+10.1875";
			elsif QstateRE(3) = to_sfixed(10.2500,QstateRE(3)) then
				char3RE <= "+10.2500";
			elsif QstateRE(3) = to_sfixed(10.3125,QstateRE(3)) then
				char3RE <= "+10.3125";
			elsif QstateRE(3) = to_sfixed(10.3750,QstateRE(3)) then
				char3RE <= "+10.3750";
			elsif QstateRE(3) = to_sfixed(10.4375,QstateRE(3)) then
				char3RE <= "+10.4375";
			elsif QstateRE(3) = to_sfixed(10.5000,QstateRE(3)) then
				char3RE <= "+10.5000";
			elsif QstateRE(3) = to_sfixed(10.5625,QstateRE(3)) then
				char3RE <= "+10.5625";
			elsif QstateRE(3) = to_sfixed(10.6250,QstateRE(3)) then
				char3RE <= "+10.6250";
			elsif QstateRE(3) = to_sfixed(10.6875,QstateRE(3)) then
				char3RE <= "+10.6875";
			elsif QstateRE(3) = to_sfixed(10.7500,QstateRE(3)) then
				char3RE <= "+10.7500";
			elsif QstateRE(3) = to_sfixed(10.8125,QstateRE(3)) then
				char3RE <= "+10.8125";
			elsif QstateRE(3) = to_sfixed(10.8750,QstateRE(3)) then
				char3RE <= "+10.8750";
			elsif QstateRE(3) = to_sfixed(10.9375,QstateRE(3)) then
				char3RE <= "+10.9375";
			elsif QstateRE(3) = to_sfixed(11.0000,QstateRE(3)) then
				char3RE <= "+11.0000";
			elsif QstateRE(3) = to_sfixed(11.0625,QstateRE(3)) then
				char3RE <= "+11.0625";
			elsif QstateRE(3) = to_sfixed(11.1250,QstateRE(3)) then
				char3RE <= "+11.1250";
			elsif QstateRE(3) = to_sfixed(11.1875,QstateRE(3)) then
				char3RE <= "+11.1875";
			elsif QstateRE(3) = to_sfixed(11.2500,QstateRE(3)) then
				char3RE <= "+11.2500";
			elsif QstateRE(3) = to_sfixed(11.3125,QstateRE(3)) then
				char3RE <= "+11.3125";
			elsif QstateRE(3) = to_sfixed(11.3750,QstateRE(3)) then
				char3RE <= "+11.3750";
			elsif QstateRE(3) = to_sfixed(11.4375,QstateRE(3)) then
				char3RE <= "+11.4375";
			elsif QstateRE(3) = to_sfixed(11.5000,QstateRE(3)) then
				char3RE <= "+11.5000";
			elsif QstateRE(3) = to_sfixed(11.5625,QstateRE(3)) then
				char3RE <= "+11.5625";
			elsif QstateRE(3) = to_sfixed(11.6250,QstateRE(3)) then
				char3RE <= "+11.6250";
			elsif QstateRE(3) = to_sfixed(11.6875,QstateRE(3)) then
				char3RE <= "+11.6875";
			elsif QstateRE(3) = to_sfixed(11.7500,QstateRE(3)) then
				char3RE <= "+11.7500";
			elsif QstateRE(3) = to_sfixed(11.8125,QstateRE(3)) then
				char3RE <= "+11.8125";
			elsif QstateRE(3) = to_sfixed(11.8750,QstateRE(3)) then
				char3RE <= "+11.8750";
			elsif QstateRE(3) = to_sfixed(11.9375,QstateRE(3)) then
				char3RE <= "+11.9375";
			elsif QstateRE(3) = to_sfixed(12.0000,QstateRE(3)) then
				char3RE <= "+12.0000";
			elsif QstateRE(3) = to_sfixed(12.0625,QstateRE(3)) then
				char3RE <= "+12.0625";
			elsif QstateRE(3) = to_sfixed(12.1250,QstateRE(3)) then
				char3RE <= "+12.1250";
			elsif QstateRE(3) = to_sfixed(12.1875,QstateRE(3)) then
				char3RE <= "+12.1875";
			elsif QstateRE(3) = to_sfixed(12.2500,QstateRE(3)) then
				char3RE <= "+12.2500";
			elsif QstateRE(3) = to_sfixed(12.3125,QstateRE(3)) then
				char3RE <= "+12.3125";
			elsif QstateRE(3) = to_sfixed(12.3750,QstateRE(3)) then
				char3RE <= "+12.3750";
			elsif QstateRE(3) = to_sfixed(12.4375,QstateRE(3)) then
				char3RE <= "+12.4375";
			elsif QstateRE(3) = to_sfixed(12.5000,QstateRE(3)) then
				char3RE <= "+12.5000";
			elsif QstateRE(3) = to_sfixed(12.5625,QstateRE(3)) then
				char3RE <= "+12.5625";
			elsif QstateRE(3) = to_sfixed(12.6250,QstateRE(3)) then
				char3RE <= "+12.6250";
			elsif QstateRE(3) = to_sfixed(12.6875,QstateRE(3)) then
				char3RE <= "+12.6875";
			elsif QstateRE(3) = to_sfixed(12.7500,QstateRE(3)) then
				char3RE <= "+12.7500";
			elsif QstateRE(3) = to_sfixed(12.8125,QstateRE(3)) then
				char3RE <= "+12.8125";
			elsif QstateRE(3) = to_sfixed(12.8750,QstateRE(3)) then
				char3RE <= "+12.8750";
			elsif QstateRE(3) = to_sfixed(12.9375,QstateRE(3)) then
				char3RE <= "+12.9375";
			elsif QstateRE(3) = to_sfixed(13.0000,QstateRE(3)) then
				char3RE <= "+13.0000";
			elsif QstateRE(3) = to_sfixed(13.0625,QstateRE(3)) then
				char3RE <= "+13.0625";
			elsif QstateRE(3) = to_sfixed(13.1250,QstateRE(3)) then
				char3RE <= "+13.1250";
			elsif QstateRE(3) = to_sfixed(13.1875,QstateRE(3)) then
				char3RE <= "+13.1875";
			elsif QstateRE(3) = to_sfixed(13.2500,QstateRE(3)) then
				char3RE <= "+13.2500";
			elsif QstateRE(3) = to_sfixed(13.3125,QstateRE(3)) then
				char3RE <= "+13.3125";
			elsif QstateRE(3) = to_sfixed(13.3750,QstateRE(3)) then
				char3RE <= "+13.3750";
			elsif QstateRE(3) = to_sfixed(13.4375,QstateRE(3)) then
				char3RE <= "+13.4375";
			elsif QstateRE(3) = to_sfixed(13.5000,QstateRE(3)) then
				char3RE <= "+13.5000";
			elsif QstateRE(3) = to_sfixed(13.5625,QstateRE(3)) then
				char3RE <= "+13.5625";
			elsif QstateRE(3) = to_sfixed(13.6250,QstateRE(3)) then
				char3RE <= "+13.6250";
			elsif QstateRE(3) = to_sfixed(13.6875,QstateRE(3)) then
				char3RE <= "+13.6875";
			elsif QstateRE(3) = to_sfixed(13.7500,QstateRE(3)) then
				char3RE <= "+13.7500";
			elsif QstateRE(3) = to_sfixed(13.8125,QstateRE(3)) then
				char3RE <= "+13.8125";
			elsif QstateRE(3) = to_sfixed(13.8750,QstateRE(3)) then
				char3RE <= "+13.8750";
			elsif QstateRE(3) = to_sfixed(13.9375,QstateRE(3)) then
				char3RE <= "+13.9375";
			elsif QstateRE(3) = to_sfixed(14.0000,QstateRE(3)) then
				char3RE <= "+14.0000";
			elsif QstateRE(3) = to_sfixed(14.0625,QstateRE(3)) then
				char3RE <= "+14.0625";
			elsif QstateRE(3) = to_sfixed(14.1250,QstateRE(3)) then
				char3RE <= "+14.1250";
			elsif QstateRE(3) = to_sfixed(14.1875,QstateRE(3)) then
				char3RE <= "+14.1875";
			elsif QstateRE(3) = to_sfixed(14.2500,QstateRE(3)) then
				char3RE <= "+14.2500";
			elsif QstateRE(3) = to_sfixed(14.3125,QstateRE(3)) then
				char3RE <= "+14.3125";
			elsif QstateRE(3) = to_sfixed(14.3750,QstateRE(3)) then
				char3RE <= "+14.3750";
			elsif QstateRE(3) = to_sfixed(14.4375,QstateRE(3)) then
				char3RE <= "+14.4375";
			elsif QstateRE(3) = to_sfixed(14.5000,QstateRE(3)) then
				char3RE <= "+14.5000";
			elsif QstateRE(3) = to_sfixed(14.5625,QstateRE(3)) then
				char3RE <= "+14.5625";
			elsif QstateRE(3) = to_sfixed(14.6250,QstateRE(3)) then
				char3RE <= "+14.6250";
			elsif QstateRE(3) = to_sfixed(14.6875,QstateRE(3)) then
				char3RE <= "+14.6875";
			elsif QstateRE(3) = to_sfixed(14.7500,QstateRE(3)) then
				char3RE <= "+14.7500";
			elsif QstateRE(3) = to_sfixed(14.8125,QstateRE(3)) then
				char3RE <= "+14.8125";
			elsif QstateRE(3) = to_sfixed(14.8750,QstateRE(3)) then
				char3RE <= "+14.8750";
			elsif QstateRE(3) = to_sfixed(14.9375,QstateRE(3)) then
				char3RE <= "+14.9375";
			elsif QstateRE(3) = to_sfixed(15.0000,QstateRE(3)) then
				char3RE <= "+15.0000";
			elsif QstateRE(3) = to_sfixed(15.0625,QstateRE(3)) then
				char3RE <= "+15.0625";
			elsif QstateRE(3) = to_sfixed(15.1250,QstateRE(3)) then
				char3RE <= "+15.1250";
			elsif QstateRE(3) = to_sfixed(15.1875,QstateRE(3)) then
				char3RE <= "+15.1875";
			elsif QstateRE(3) = to_sfixed(15.2500,QstateRE(3)) then
				char3RE <= "+15.2500";
			elsif QstateRE(3) = to_sfixed(15.3125,QstateRE(3)) then
				char3RE <= "+15.3125";
			elsif QstateRE(3) = to_sfixed(15.3750,QstateRE(3)) then
				char3RE <= "+15.3750";
			elsif QstateRE(3) = to_sfixed(15.4375,QstateRE(3)) then
				char3RE <= "+15.4375";
			elsif QstateRE(3) = to_sfixed(15.5000,QstateRE(3)) then
				char3RE <= "+15.5000";
			elsif QstateRE(3) = to_sfixed(15.5625,QstateRE(3)) then
				char3RE <= "+15.5625";
			elsif QstateRE(3) = to_sfixed(15.6250,QstateRE(3)) then
				char3RE <= "+15.6250";
			elsif QstateRE(3) = to_sfixed(15.6875,QstateRE(3)) then
				char3RE <= "+15.6875";
			elsif QstateRE(3) = to_sfixed(15.7500,QstateRE(3)) then
				char3RE <= "+15.7500";
			elsif QstateRE(3) = to_sfixed(15.8125,QstateRE(3)) then
				char3RE <= "+15.8125";
			elsif QstateRE(3) = to_sfixed(15.8750,QstateRE(3)) then
				char3RE <= "+15.8750";
			elsif QstateRE(3) = to_sfixed(15.9375,QstateRE(3)) then
				char3RE <= "+15.9375";
			end if;
			if QstateIM(3) = to_sfixed(-15.9375,QstateIM(3)) then
				char3IM <= "-15.9375";
			elsif QstateIM(3) = to_sfixed(-15.8750,QstateIM(3)) then
				char3IM <= "-15.8750";
			elsif QstateIM(3) = to_sfixed(-15.8125,QstateIM(3)) then
				char3IM <= "-15.8125";
			elsif QstateIM(3) = to_sfixed(-15.7500,QstateIM(3)) then
				char3IM <= "-15.7500";
			elsif QstateIM(3) = to_sfixed(-15.6875,QstateIM(3)) then
				char3IM <= "-15.6875";
			elsif QstateIM(3) = to_sfixed(-15.6250,QstateIM(3)) then
				char3IM <= "-15.6250";
			elsif QstateIM(3) = to_sfixed(-15.5625,QstateIM(3)) then
				char3IM <= "-15.5625";
			elsif QstateIM(3) = to_sfixed(-15.5000,QstateIM(3)) then
				char3IM <= "-15.5000";
			elsif QstateIM(3) = to_sfixed(-15.4375,QstateIM(3)) then
				char3IM <= "-15.4375";
			elsif QstateIM(3) = to_sfixed(-15.3750,QstateIM(3)) then
				char3IM <= "-15.3750";
			elsif QstateIM(3) = to_sfixed(-15.3125,QstateIM(3)) then
				char3IM <= "-15.3125";
			elsif QstateIM(3) = to_sfixed(-15.2500,QstateIM(3)) then
				char3IM <= "-15.2500";
			elsif QstateIM(3) = to_sfixed(-15.1875,QstateIM(3)) then
				char3IM <= "-15.1875";
			elsif QstateIM(3) = to_sfixed(-15.1250,QstateIM(3)) then
				char3IM <= "-15.1250";
			elsif QstateIM(3) = to_sfixed(-15.0625,QstateIM(3)) then
				char3IM <= "-15.0625";
			elsif QstateIM(3) = to_sfixed(-15.0000,QstateIM(3)) then
				char3IM <= "-15.0000";
			elsif QstateIM(3) = to_sfixed(-14.9375,QstateIM(3)) then
				char3IM <= "-14.9375";
			elsif QstateIM(3) = to_sfixed(-14.8750,QstateIM(3)) then
				char3IM <= "-14.8750";
			elsif QstateIM(3) = to_sfixed(-14.8125,QstateIM(3)) then
				char3IM <= "-14.8125";
			elsif QstateIM(3) = to_sfixed(-14.7500,QstateIM(3)) then
				char3IM <= "-14.7500";
			elsif QstateIM(3) = to_sfixed(-14.6875,QstateIM(3)) then
				char3IM <= "-14.6875";
			elsif QstateIM(3) = to_sfixed(-14.6250,QstateIM(3)) then
				char3IM <= "-14.6250";
			elsif QstateIM(3) = to_sfixed(-14.5625,QstateIM(3)) then
				char3IM <= "-14.5625";
			elsif QstateIM(3) = to_sfixed(-14.5000,QstateIM(3)) then
				char3IM <= "-14.5000";
			elsif QstateIM(3) = to_sfixed(-14.4375,QstateIM(3)) then
				char3IM <= "-14.4375";
			elsif QstateIM(3) = to_sfixed(-14.3750,QstateIM(3)) then
				char3IM <= "-14.3750";
			elsif QstateIM(3) = to_sfixed(-14.3125,QstateIM(3)) then
				char3IM <= "-14.3125";
			elsif QstateIM(3) = to_sfixed(-14.2500,QstateIM(3)) then
				char3IM <= "-14.2500";
			elsif QstateIM(3) = to_sfixed(-14.1875,QstateIM(3)) then
				char3IM <= "-14.1875";
			elsif QstateIM(3) = to_sfixed(-14.1250,QstateIM(3)) then
				char3IM <= "-14.1250";
			elsif QstateIM(3) = to_sfixed(-14.0625,QstateIM(3)) then
				char3IM <= "-14.0625";
			elsif QstateIM(3) = to_sfixed(-14.0000,QstateIM(3)) then
				char3IM <= "-14.0000";
			elsif QstateIM(3) = to_sfixed(-13.9375,QstateIM(3)) then
				char3IM <= "-13.9375";
			elsif QstateIM(3) = to_sfixed(-13.8750,QstateIM(3)) then
				char3IM <= "-13.8750";
			elsif QstateIM(3) = to_sfixed(-13.8125,QstateIM(3)) then
				char3IM <= "-13.8125";
			elsif QstateIM(3) = to_sfixed(-13.7500,QstateIM(3)) then
				char3IM <= "-13.7500";
			elsif QstateIM(3) = to_sfixed(-13.6875,QstateIM(3)) then
				char3IM <= "-13.6875";
			elsif QstateIM(3) = to_sfixed(-13.6250,QstateIM(3)) then
				char3IM <= "-13.6250";
			elsif QstateIM(3) = to_sfixed(-13.5625,QstateIM(3)) then
				char3IM <= "-13.5625";
			elsif QstateIM(3) = to_sfixed(-13.5000,QstateIM(3)) then
				char3IM <= "-13.5000";
			elsif QstateIM(3) = to_sfixed(-13.4375,QstateIM(3)) then
				char3IM <= "-13.4375";
			elsif QstateIM(3) = to_sfixed(-13.3750,QstateIM(3)) then
				char3IM <= "-13.3750";
			elsif QstateIM(3) = to_sfixed(-13.3125,QstateIM(3)) then
				char3IM <= "-13.3125";
			elsif QstateIM(3) = to_sfixed(-13.2500,QstateIM(3)) then
				char3IM <= "-13.2500";
			elsif QstateIM(3) = to_sfixed(-13.1875,QstateIM(3)) then
				char3IM <= "-13.1875";
			elsif QstateIM(3) = to_sfixed(-13.1250,QstateIM(3)) then
				char3IM <= "-13.1250";
			elsif QstateIM(3) = to_sfixed(-13.0625,QstateIM(3)) then
				char3IM <= "-13.0625";
			elsif QstateIM(3) = to_sfixed(-13.0000,QstateIM(3)) then
				char3IM <= "-13.0000";
			elsif QstateIM(3) = to_sfixed(-12.9375,QstateIM(3)) then
				char3IM <= "-12.9375";
			elsif QstateIM(3) = to_sfixed(-12.8750,QstateIM(3)) then
				char3IM <= "-12.8750";
			elsif QstateIM(3) = to_sfixed(-12.8125,QstateIM(3)) then
				char3IM <= "-12.8125";
			elsif QstateIM(3) = to_sfixed(-12.7500,QstateIM(3)) then
				char3IM <= "-12.7500";
			elsif QstateIM(3) = to_sfixed(-12.6875,QstateIM(3)) then
				char3IM <= "-12.6875";
			elsif QstateIM(3) = to_sfixed(-12.6250,QstateIM(3)) then
				char3IM <= "-12.6250";
			elsif QstateIM(3) = to_sfixed(-12.5625,QstateIM(3)) then
				char3IM <= "-12.5625";
			elsif QstateIM(3) = to_sfixed(-12.5000,QstateIM(3)) then
				char3IM <= "-12.5000";
			elsif QstateIM(3) = to_sfixed(-12.4375,QstateIM(3)) then
				char3IM <= "-12.4375";
			elsif QstateIM(3) = to_sfixed(-12.3750,QstateIM(3)) then
				char3IM <= "-12.3750";
			elsif QstateIM(3) = to_sfixed(-12.3125,QstateIM(3)) then
				char3IM <= "-12.3125";
			elsif QstateIM(3) = to_sfixed(-12.2500,QstateIM(3)) then
				char3IM <= "-12.2500";
			elsif QstateIM(3) = to_sfixed(-12.1875,QstateIM(3)) then
				char3IM <= "-12.1875";
			elsif QstateIM(3) = to_sfixed(-12.1250,QstateIM(3)) then
				char3IM <= "-12.1250";
			elsif QstateIM(3) = to_sfixed(-12.0625,QstateIM(3)) then
				char3IM <= "-12.0625";
			elsif QstateIM(3) = to_sfixed(-12.0000,QstateIM(3)) then
				char3IM <= "-12.0000";
			elsif QstateIM(3) = to_sfixed(-11.9375,QstateIM(3)) then
				char3IM <= "-11.9375";
			elsif QstateIM(3) = to_sfixed(-11.8750,QstateIM(3)) then
				char3IM <= "-11.8750";
			elsif QstateIM(3) = to_sfixed(-11.8125,QstateIM(3)) then
				char3IM <= "-11.8125";
			elsif QstateIM(3) = to_sfixed(-11.7500,QstateIM(3)) then
				char3IM <= "-11.7500";
			elsif QstateIM(3) = to_sfixed(-11.6875,QstateIM(3)) then
				char3IM <= "-11.6875";
			elsif QstateIM(3) = to_sfixed(-11.6250,QstateIM(3)) then
				char3IM <= "-11.6250";
			elsif QstateIM(3) = to_sfixed(-11.5625,QstateIM(3)) then
				char3IM <= "-11.5625";
			elsif QstateIM(3) = to_sfixed(-11.5000,QstateIM(3)) then
				char3IM <= "-11.5000";
			elsif QstateIM(3) = to_sfixed(-11.4375,QstateIM(3)) then
				char3IM <= "-11.4375";
			elsif QstateIM(3) = to_sfixed(-11.3750,QstateIM(3)) then
				char3IM <= "-11.3750";
			elsif QstateIM(3) = to_sfixed(-11.3125,QstateIM(3)) then
				char3IM <= "-11.3125";
			elsif QstateIM(3) = to_sfixed(-11.2500,QstateIM(3)) then
				char3IM <= "-11.2500";
			elsif QstateIM(3) = to_sfixed(-11.1875,QstateIM(3)) then
				char3IM <= "-11.1875";
			elsif QstateIM(3) = to_sfixed(-11.1250,QstateIM(3)) then
				char3IM <= "-11.1250";
			elsif QstateIM(3) = to_sfixed(-11.0625,QstateIM(3)) then
				char3IM <= "-11.0625";
			elsif QstateIM(3) = to_sfixed(-11.0000,QstateIM(3)) then
				char3IM <= "-11.0000";
			elsif QstateIM(3) = to_sfixed(-10.9375,QstateIM(3)) then
				char3IM <= "-10.9375";
			elsif QstateIM(3) = to_sfixed(-10.8750,QstateIM(3)) then
				char3IM <= "-10.8750";
			elsif QstateIM(3) = to_sfixed(-10.8125,QstateIM(3)) then
				char3IM <= "-10.8125";
			elsif QstateIM(3) = to_sfixed(-10.7500,QstateIM(3)) then
				char3IM <= "-10.7500";
			elsif QstateIM(3) = to_sfixed(-10.6875,QstateIM(3)) then
				char3IM <= "-10.6875";
			elsif QstateIM(3) = to_sfixed(-10.6250,QstateIM(3)) then
				char3IM <= "-10.6250";
			elsif QstateIM(3) = to_sfixed(-10.5625,QstateIM(3)) then
				char3IM <= "-10.5625";
			elsif QstateIM(3) = to_sfixed(-10.5000,QstateIM(3)) then
				char3IM <= "-10.5000";
			elsif QstateIM(3) = to_sfixed(-10.4375,QstateIM(3)) then
				char3IM <= "-10.4375";
			elsif QstateIM(3) = to_sfixed(-10.3750,QstateIM(3)) then
				char3IM <= "-10.3750";
			elsif QstateIM(3) = to_sfixed(-10.3125,QstateIM(3)) then
				char3IM <= "-10.3125";
			elsif QstateIM(3) = to_sfixed(-10.2500,QstateIM(3)) then
				char3IM <= "-10.2500";
			elsif QstateIM(3) = to_sfixed(-10.1875,QstateIM(3)) then
				char3IM <= "-10.1875";
			elsif QstateIM(3) = to_sfixed(-10.1250,QstateIM(3)) then
				char3IM <= "-10.1250";
			elsif QstateIM(3) = to_sfixed(-10.0625,QstateIM(3)) then
				char3IM <= "-10.0625";
			elsif QstateIM(3) = to_sfixed(-10.0000,QstateIM(3)) then
				char3IM <= "-10.0000";
			elsif QstateIM(3) = to_sfixed(-9.9375,QstateIM(3)) then
				char3IM <= "--9.9375";
			elsif QstateIM(3) = to_sfixed(-9.8750,QstateIM(3)) then
				char3IM <= "--9.8750";
			elsif QstateIM(3) = to_sfixed(-9.8125,QstateIM(3)) then
				char3IM <= "--9.8125";
			elsif QstateIM(3) = to_sfixed(-9.7500,QstateIM(3)) then
				char3IM <= "--9.7500";
			elsif QstateIM(3) = to_sfixed(-9.6875,QstateIM(3)) then
				char3IM <= "--9.6875";
			elsif QstateIM(3) = to_sfixed(-9.6250,QstateIM(3)) then
				char3IM <= "--9.6250";
			elsif QstateIM(3) = to_sfixed(-9.5625,QstateIM(3)) then
				char3IM <= "--9.5625";
			elsif QstateIM(3) = to_sfixed(-9.5000,QstateIM(3)) then
				char3IM <= "--9.5000";
			elsif QstateIM(3) = to_sfixed(-9.4375,QstateIM(3)) then
				char3IM <= "--9.4375";
			elsif QstateIM(3) = to_sfixed(-9.3750,QstateIM(3)) then
				char3IM <= "--9.3750";
			elsif QstateIM(3) = to_sfixed(-9.3125,QstateIM(3)) then
				char3IM <= "--9.3125";
			elsif QstateIM(3) = to_sfixed(-9.2500,QstateIM(3)) then
				char3IM <= "--9.2500";
			elsif QstateIM(3) = to_sfixed(-9.1875,QstateIM(3)) then
				char3IM <= "--9.1875";
			elsif QstateIM(3) = to_sfixed(-9.1250,QstateIM(3)) then
				char3IM <= "--9.1250";
			elsif QstateIM(3) = to_sfixed(-9.0625,QstateIM(3)) then
				char3IM <= "--9.0625";
			elsif QstateIM(3) = to_sfixed(-9.0000,QstateIM(3)) then
				char3IM <= "--9.0000";
			elsif QstateIM(3) = to_sfixed(-8.9375,QstateIM(3)) then
				char3IM <= "--8.9375";
			elsif QstateIM(3) = to_sfixed(-8.8750,QstateIM(3)) then
				char3IM <= "--8.8750";
			elsif QstateIM(3) = to_sfixed(-8.8125,QstateIM(3)) then
				char3IM <= "--8.8125";
			elsif QstateIM(3) = to_sfixed(-8.7500,QstateIM(3)) then
				char3IM <= "--8.7500";
			elsif QstateIM(3) = to_sfixed(-8.6875,QstateIM(3)) then
				char3IM <= "--8.6875";
			elsif QstateIM(3) = to_sfixed(-8.6250,QstateIM(3)) then
				char3IM <= "--8.6250";
			elsif QstateIM(3) = to_sfixed(-8.5625,QstateIM(3)) then
				char3IM <= "--8.5625";
			elsif QstateIM(3) = to_sfixed(-8.5000,QstateIM(3)) then
				char3IM <= "--8.5000";
			elsif QstateIM(3) = to_sfixed(-8.4375,QstateIM(3)) then
				char3IM <= "--8.4375";
			elsif QstateIM(3) = to_sfixed(-8.3750,QstateIM(3)) then
				char3IM <= "--8.3750";
			elsif QstateIM(3) = to_sfixed(-8.3125,QstateIM(3)) then
				char3IM <= "--8.3125";
			elsif QstateIM(3) = to_sfixed(-8.2500,QstateIM(3)) then
				char3IM <= "--8.2500";
			elsif QstateIM(3) = to_sfixed(-8.1875,QstateIM(3)) then
				char3IM <= "--8.1875";
			elsif QstateIM(3) = to_sfixed(-8.1250,QstateIM(3)) then
				char3IM <= "--8.1250";
			elsif QstateIM(3) = to_sfixed(-8.0625,QstateIM(3)) then
				char3IM <= "--8.0625";
			elsif QstateIM(3) = to_sfixed(-8.0000,QstateIM(3)) then
				char3IM <= "--8.0000";
			elsif QstateIM(3) = to_sfixed(-7.9375,QstateIM(3)) then
				char3IM <= "--7.9375";
			elsif QstateIM(3) = to_sfixed(-7.8750,QstateIM(3)) then
				char3IM <= "--7.8750";
			elsif QstateIM(3) = to_sfixed(-7.8125,QstateIM(3)) then
				char3IM <= "--7.8125";
			elsif QstateIM(3) = to_sfixed(-7.7500,QstateIM(3)) then
				char3IM <= "--7.7500";
			elsif QstateIM(3) = to_sfixed(-7.6875,QstateIM(3)) then
				char3IM <= "--7.6875";
			elsif QstateIM(3) = to_sfixed(-7.6250,QstateIM(3)) then
				char3IM <= "--7.6250";
			elsif QstateIM(3) = to_sfixed(-7.5625,QstateIM(3)) then
				char3IM <= "--7.5625";
			elsif QstateIM(3) = to_sfixed(-7.5000,QstateIM(3)) then
				char3IM <= "--7.5000";
			elsif QstateIM(3) = to_sfixed(-7.4375,QstateIM(3)) then
				char3IM <= "--7.4375";
			elsif QstateIM(3) = to_sfixed(-7.3750,QstateIM(3)) then
				char3IM <= "--7.3750";
			elsif QstateIM(3) = to_sfixed(-7.3125,QstateIM(3)) then
				char3IM <= "--7.3125";
			elsif QstateIM(3) = to_sfixed(-7.2500,QstateIM(3)) then
				char3IM <= "--7.2500";
			elsif QstateIM(3) = to_sfixed(-7.1875,QstateIM(3)) then
				char3IM <= "--7.1875";
			elsif QstateIM(3) = to_sfixed(-7.1250,QstateIM(3)) then
				char3IM <= "--7.1250";
			elsif QstateIM(3) = to_sfixed(-7.0625,QstateIM(3)) then
				char3IM <= "--7.0625";
			elsif QstateIM(3) = to_sfixed(-7.0000,QstateIM(3)) then
				char3IM <= "--7.0000";
			elsif QstateIM(3) = to_sfixed(-6.9375,QstateIM(3)) then
				char3IM <= "--6.9375";
			elsif QstateIM(3) = to_sfixed(-6.8750,QstateIM(3)) then
				char3IM <= "--6.8750";
			elsif QstateIM(3) = to_sfixed(-6.8125,QstateIM(3)) then
				char3IM <= "--6.8125";
			elsif QstateIM(3) = to_sfixed(-6.7500,QstateIM(3)) then
				char3IM <= "--6.7500";
			elsif QstateIM(3) = to_sfixed(-6.6875,QstateIM(3)) then
				char3IM <= "--6.6875";
			elsif QstateIM(3) = to_sfixed(-6.6250,QstateIM(3)) then
				char3IM <= "--6.6250";
			elsif QstateIM(3) = to_sfixed(-6.5625,QstateIM(3)) then
				char3IM <= "--6.5625";
			elsif QstateIM(3) = to_sfixed(-6.5000,QstateIM(3)) then
				char3IM <= "--6.5000";
			elsif QstateIM(3) = to_sfixed(-6.4375,QstateIM(3)) then
				char3IM <= "--6.4375";
			elsif QstateIM(3) = to_sfixed(-6.3750,QstateIM(3)) then
				char3IM <= "--6.3750";
			elsif QstateIM(3) = to_sfixed(-6.3125,QstateIM(3)) then
				char3IM <= "--6.3125";
			elsif QstateIM(3) = to_sfixed(-6.2500,QstateIM(3)) then
				char3IM <= "--6.2500";
			elsif QstateIM(3) = to_sfixed(-6.1875,QstateIM(3)) then
				char3IM <= "--6.1875";
			elsif QstateIM(3) = to_sfixed(-6.1250,QstateIM(3)) then
				char3IM <= "--6.1250";
			elsif QstateIM(3) = to_sfixed(-6.0625,QstateIM(3)) then
				char3IM <= "--6.0625";
			elsif QstateIM(3) = to_sfixed(-6.0000,QstateIM(3)) then
				char3IM <= "--6.0000";
			elsif QstateIM(3) = to_sfixed(-5.9375,QstateIM(3)) then
				char3IM <= "--5.9375";
			elsif QstateIM(3) = to_sfixed(-5.8750,QstateIM(3)) then
				char3IM <= "--5.8750";
			elsif QstateIM(3) = to_sfixed(-5.8125,QstateIM(3)) then
				char3IM <= "--5.8125";
			elsif QstateIM(3) = to_sfixed(-5.7500,QstateIM(3)) then
				char3IM <= "--5.7500";
			elsif QstateIM(3) = to_sfixed(-5.6875,QstateIM(3)) then
				char3IM <= "--5.6875";
			elsif QstateIM(3) = to_sfixed(-5.6250,QstateIM(3)) then
				char3IM <= "--5.6250";
			elsif QstateIM(3) = to_sfixed(-5.5625,QstateIM(3)) then
				char3IM <= "--5.5625";
			elsif QstateIM(3) = to_sfixed(-5.5000,QstateIM(3)) then
				char3IM <= "--5.5000";
			elsif QstateIM(3) = to_sfixed(-5.4375,QstateIM(3)) then
				char3IM <= "--5.4375";
			elsif QstateIM(3) = to_sfixed(-5.3750,QstateIM(3)) then
				char3IM <= "--5.3750";
			elsif QstateIM(3) = to_sfixed(-5.3125,QstateIM(3)) then
				char3IM <= "--5.3125";
			elsif QstateIM(3) = to_sfixed(-5.2500,QstateIM(3)) then
				char3IM <= "--5.2500";
			elsif QstateIM(3) = to_sfixed(-5.1875,QstateIM(3)) then
				char3IM <= "--5.1875";
			elsif QstateIM(3) = to_sfixed(-5.1250,QstateIM(3)) then
				char3IM <= "--5.1250";
			elsif QstateIM(3) = to_sfixed(-5.0625,QstateIM(3)) then
				char3IM <= "--5.0625";
			elsif QstateIM(3) = to_sfixed(-5.0000,QstateIM(3)) then
				char3IM <= "--5.0000";
			elsif QstateIM(3) = to_sfixed(-4.9375,QstateIM(3)) then
				char3IM <= "--4.9375";
			elsif QstateIM(3) = to_sfixed(-4.8750,QstateIM(3)) then
				char3IM <= "--4.8750";
			elsif QstateIM(3) = to_sfixed(-4.8125,QstateIM(3)) then
				char3IM <= "--4.8125";
			elsif QstateIM(3) = to_sfixed(-4.7500,QstateIM(3)) then
				char3IM <= "--4.7500";
			elsif QstateIM(3) = to_sfixed(-4.6875,QstateIM(3)) then
				char3IM <= "--4.6875";
			elsif QstateIM(3) = to_sfixed(-4.6250,QstateIM(3)) then
				char3IM <= "--4.6250";
			elsif QstateIM(3) = to_sfixed(-4.5625,QstateIM(3)) then
				char3IM <= "--4.5625";
			elsif QstateIM(3) = to_sfixed(-4.5000,QstateIM(3)) then
				char3IM <= "--4.5000";
			elsif QstateIM(3) = to_sfixed(-4.4375,QstateIM(3)) then
				char3IM <= "--4.4375";
			elsif QstateIM(3) = to_sfixed(-4.3750,QstateIM(3)) then
				char3IM <= "--4.3750";
			elsif QstateIM(3) = to_sfixed(-4.3125,QstateIM(3)) then
				char3IM <= "--4.3125";
			elsif QstateIM(3) = to_sfixed(-4.2500,QstateIM(3)) then
				char3IM <= "--4.2500";
			elsif QstateIM(3) = to_sfixed(-4.1875,QstateIM(3)) then
				char3IM <= "--4.1875";
			elsif QstateIM(3) = to_sfixed(-4.1250,QstateIM(3)) then
				char3IM <= "--4.1250";
			elsif QstateIM(3) = to_sfixed(-4.0625,QstateIM(3)) then
				char3IM <= "--4.0625";
			elsif QstateIM(3) = to_sfixed(-4.0000,QstateIM(3)) then
				char3IM <= "--4.0000";
			elsif QstateIM(3) = to_sfixed(-3.9375,QstateIM(3)) then
				char3IM <= "--3.9375";
			elsif QstateIM(3) = to_sfixed(-3.8750,QstateIM(3)) then
				char3IM <= "--3.8750";
			elsif QstateIM(3) = to_sfixed(-3.8125,QstateIM(3)) then
				char3IM <= "--3.8125";
			elsif QstateIM(3) = to_sfixed(-3.7500,QstateIM(3)) then
				char3IM <= "--3.7500";
			elsif QstateIM(3) = to_sfixed(-3.6875,QstateIM(3)) then
				char3IM <= "--3.6875";
			elsif QstateIM(3) = to_sfixed(-3.6250,QstateIM(3)) then
				char3IM <= "--3.6250";
			elsif QstateIM(3) = to_sfixed(-3.5625,QstateIM(3)) then
				char3IM <= "--3.5625";
			elsif QstateIM(3) = to_sfixed(-3.5000,QstateIM(3)) then
				char3IM <= "--3.5000";
			elsif QstateIM(3) = to_sfixed(-3.4375,QstateIM(3)) then
				char3IM <= "--3.4375";
			elsif QstateIM(3) = to_sfixed(-3.3750,QstateIM(3)) then
				char3IM <= "--3.3750";
			elsif QstateIM(3) = to_sfixed(-3.3125,QstateIM(3)) then
				char3IM <= "--3.3125";
			elsif QstateIM(3) = to_sfixed(-3.2500,QstateIM(3)) then
				char3IM <= "--3.2500";
			elsif QstateIM(3) = to_sfixed(-3.1875,QstateIM(3)) then
				char3IM <= "--3.1875";
			elsif QstateIM(3) = to_sfixed(-3.1250,QstateIM(3)) then
				char3IM <= "--3.1250";
			elsif QstateIM(3) = to_sfixed(-3.0625,QstateIM(3)) then
				char3IM <= "--3.0625";
			elsif QstateIM(3) = to_sfixed(-3.0000,QstateIM(3)) then
				char3IM <= "--3.0000";
			elsif QstateIM(3) = to_sfixed(-2.9375,QstateIM(3)) then
				char3IM <= "--2.9375";
			elsif QstateIM(3) = to_sfixed(-2.8750,QstateIM(3)) then
				char3IM <= "--2.8750";
			elsif QstateIM(3) = to_sfixed(-2.8125,QstateIM(3)) then
				char3IM <= "--2.8125";
			elsif QstateIM(3) = to_sfixed(-2.7500,QstateIM(3)) then
				char3IM <= "--2.7500";
			elsif QstateIM(3) = to_sfixed(-2.6875,QstateIM(3)) then
				char3IM <= "--2.6875";
			elsif QstateIM(3) = to_sfixed(-2.6250,QstateIM(3)) then
				char3IM <= "--2.6250";
			elsif QstateIM(3) = to_sfixed(-2.5625,QstateIM(3)) then
				char3IM <= "--2.5625";
			elsif QstateIM(3) = to_sfixed(-2.5000,QstateIM(3)) then
				char3IM <= "--2.5000";
			elsif QstateIM(3) = to_sfixed(-2.4375,QstateIM(3)) then
				char3IM <= "--2.4375";
			elsif QstateIM(3) = to_sfixed(-2.3750,QstateIM(3)) then
				char3IM <= "--2.3750";
			elsif QstateIM(3) = to_sfixed(-2.3125,QstateIM(3)) then
				char3IM <= "--2.3125";
			elsif QstateIM(3) = to_sfixed(-2.2500,QstateIM(3)) then
				char3IM <= "--2.2500";
			elsif QstateIM(3) = to_sfixed(-2.1875,QstateIM(3)) then
				char3IM <= "--2.1875";
			elsif QstateIM(3) = to_sfixed(-2.1250,QstateIM(3)) then
				char3IM <= "--2.1250";
			elsif QstateIM(3) = to_sfixed(-2.0625,QstateIM(3)) then
				char3IM <= "--2.0625";
			elsif QstateIM(3) = to_sfixed(-2.0000,QstateIM(3)) then
				char3IM <= "--2.0000";
			elsif QstateIM(3) = to_sfixed(-1.9375,QstateIM(3)) then
				char3IM <= "--1.9375";
			elsif QstateIM(3) = to_sfixed(-1.8750,QstateIM(3)) then
				char3IM <= "--1.8750";
			elsif QstateIM(3) = to_sfixed(-1.8125,QstateIM(3)) then
				char3IM <= "--1.8125";
			elsif QstateIM(3) = to_sfixed(-1.7500,QstateIM(3)) then
				char3IM <= "--1.7500";
			elsif QstateIM(3) = to_sfixed(-1.6875,QstateIM(3)) then
				char3IM <= "--1.6875";
			elsif QstateIM(3) = to_sfixed(-1.6250,QstateIM(3)) then
				char3IM <= "--1.6250";
			elsif QstateIM(3) = to_sfixed(-1.5625,QstateIM(3)) then
				char3IM <= "--1.5625";
			elsif QstateIM(3) = to_sfixed(-1.5000,QstateIM(3)) then
				char3IM <= "--1.5000";
			elsif QstateIM(3) = to_sfixed(-1.4375,QstateIM(3)) then
				char3IM <= "--1.4375";
			elsif QstateIM(3) = to_sfixed(-1.3750,QstateIM(3)) then
				char3IM <= "--1.3750";
			elsif QstateIM(3) = to_sfixed(-1.3125,QstateIM(3)) then
				char3IM <= "--1.3125";
			elsif QstateIM(3) = to_sfixed(-1.2500,QstateIM(3)) then
				char3IM <= "--1.2500";
			elsif QstateIM(3) = to_sfixed(-1.1875,QstateIM(3)) then
				char3IM <= "--1.1875";
			elsif QstateIM(3) = to_sfixed(-1.1250,QstateIM(3)) then
				char3IM <= "--1.1250";
			elsif QstateIM(3) = to_sfixed(-1.0625,QstateIM(3)) then
				char3IM <= "--1.0625";
			elsif QstateIM(3) = to_sfixed(-1.0000,QstateIM(3)) then
				char3IM <= "--1.0000";
			elsif QstateIM(3) = to_sfixed(-0.9375,QstateIM(3)) then
				char3IM <= "--0.9375";
			elsif QstateIM(3) = to_sfixed(-0.8750,QstateIM(3)) then
				char3IM <= "--0.8750";
			elsif QstateIM(3) = to_sfixed(-0.8125,QstateIM(3)) then
				char3IM <= "--0.8125";
			elsif QstateIM(3) = to_sfixed(-0.7500,QstateIM(3)) then
				char3IM <= "--0.7500";
			elsif QstateIM(3) = to_sfixed(-0.6875,QstateIM(3)) then
				char3IM <= "--0.6875";
			elsif QstateIM(3) = to_sfixed(-0.6250,QstateIM(3)) then
				char3IM <= "--0.6250";
			elsif QstateIM(3) = to_sfixed(-0.5625,QstateIM(3)) then
				char3IM <= "--0.5625";
			elsif QstateIM(3) = to_sfixed(-0.5000,QstateIM(3)) then
				char3IM <= "--0.5000";
			elsif QstateIM(3) = to_sfixed(-0.4375,QstateIM(3)) then
				char3IM <= "--0.4375";
			elsif QstateIM(3) = to_sfixed(-0.3750,QstateIM(3)) then
				char3IM <= "--0.3750";
			elsif QstateIM(3) = to_sfixed(-0.3125,QstateIM(3)) then
				char3IM <= "--0.3125";
			elsif QstateIM(3) = to_sfixed(-0.2500,QstateIM(3)) then
				char3IM <= "--0.2500";
			elsif QstateIM(3) = to_sfixed(-0.1875,QstateIM(3)) then
				char3IM <= "--0.1875";
			elsif QstateIM(3) = to_sfixed(-0.1250,QstateIM(3)) then
				char3IM <= "--0.1250";
			elsif QstateIM(3) = to_sfixed(-0.0625,QstateIM(3)) then
				char3IM <= "--0.0625";
			elsif QstateIM(3) = to_sfixed(00.0000,QstateIM(3)) then
				char3IM <= "+00.0000";
			elsif QstateIM(3) = to_sfixed(00.0625,QstateIM(3)) then
				char3IM <= "+00.0625";
			elsif QstateIM(3) = to_sfixed(00.1250,QstateIM(3)) then
				char3IM <= "+00.1250";
			elsif QstateIM(3) = to_sfixed(00.1875,QstateIM(3)) then
				char3IM <= "+00.1875";
			elsif QstateIM(3) = to_sfixed(00.2500,QstateIM(3)) then
				char3IM <= "+00.2500";
			elsif QstateIM(3) = to_sfixed(00.3125,QstateIM(3)) then
				char3IM <= "+00.3125";
			elsif QstateIM(3) = to_sfixed(00.3750,QstateIM(3)) then
				char3IM <= "+00.3750";
			elsif QstateIM(3) = to_sfixed(00.4375,QstateIM(3)) then
				char3IM <= "+00.4375";
			elsif QstateIM(3) = to_sfixed(00.5000,QstateIM(3)) then
				char3IM <= "+00.5000";
			elsif QstateIM(3) = to_sfixed(00.5625,QstateIM(3)) then
				char3IM <= "+00.5625";
			elsif QstateIM(3) = to_sfixed(00.6250,QstateIM(3)) then
				char3IM <= "+00.6250";
			elsif QstateIM(3) = to_sfixed(00.6875,QstateIM(3)) then
				char3IM <= "+00.6875";
			elsif QstateIM(3) = to_sfixed(00.7500,QstateIM(3)) then
				char3IM <= "+00.7500";
			elsif QstateIM(3) = to_sfixed(00.8125,QstateIM(3)) then
				char3IM <= "+00.8125";
			elsif QstateIM(3) = to_sfixed(00.8750,QstateIM(3)) then
				char3IM <= "+00.8750";
			elsif QstateIM(3) = to_sfixed(00.9375,QstateIM(3)) then
				char3IM <= "+00.9375";
			elsif QstateIM(3) = to_sfixed(01.0000,QstateIM(3)) then
				char3IM <= "+01.0000";
			elsif QstateIM(3) = to_sfixed(01.0625,QstateIM(3)) then
				char3IM <= "+01.0625";
			elsif QstateIM(3) = to_sfixed(01.1250,QstateIM(3)) then
				char3IM <= "+01.1250";
			elsif QstateIM(3) = to_sfixed(01.1875,QstateIM(3)) then
				char3IM <= "+01.1875";
			elsif QstateIM(3) = to_sfixed(01.2500,QstateIM(3)) then
				char3IM <= "+01.2500";
			elsif QstateIM(3) = to_sfixed(01.3125,QstateIM(3)) then
				char3IM <= "+01.3125";
			elsif QstateIM(3) = to_sfixed(01.3750,QstateIM(3)) then
				char3IM <= "+01.3750";
			elsif QstateIM(3) = to_sfixed(01.4375,QstateIM(3)) then
				char3IM <= "+01.4375";
			elsif QstateIM(3) = to_sfixed(01.5000,QstateIM(3)) then
				char3IM <= "+01.5000";
			elsif QstateIM(3) = to_sfixed(01.5625,QstateIM(3)) then
				char3IM <= "+01.5625";
			elsif QstateIM(3) = to_sfixed(01.6250,QstateIM(3)) then
				char3IM <= "+01.6250";
			elsif QstateIM(3) = to_sfixed(01.6875,QstateIM(3)) then
				char3IM <= "+01.6875";
			elsif QstateIM(3) = to_sfixed(01.7500,QstateIM(3)) then
				char3IM <= "+01.7500";
			elsif QstateIM(3) = to_sfixed(01.8125,QstateIM(3)) then
				char3IM <= "+01.8125";
			elsif QstateIM(3) = to_sfixed(01.8750,QstateIM(3)) then
				char3IM <= "+01.8750";
			elsif QstateIM(3) = to_sfixed(01.9375,QstateIM(3)) then
				char3IM <= "+01.9375";
			elsif QstateIM(3) = to_sfixed(02.0000,QstateIM(3)) then
				char3IM <= "+02.0000";
			elsif QstateIM(3) = to_sfixed(02.0625,QstateIM(3)) then
				char3IM <= "+02.0625";
			elsif QstateIM(3) = to_sfixed(02.1250,QstateIM(3)) then
				char3IM <= "+02.1250";
			elsif QstateIM(3) = to_sfixed(02.1875,QstateIM(3)) then
				char3IM <= "+02.1875";
			elsif QstateIM(3) = to_sfixed(02.2500,QstateIM(3)) then
				char3IM <= "+02.2500";
			elsif QstateIM(3) = to_sfixed(02.3125,QstateIM(3)) then
				char3IM <= "+02.3125";
			elsif QstateIM(3) = to_sfixed(02.3750,QstateIM(3)) then
				char3IM <= "+02.3750";
			elsif QstateIM(3) = to_sfixed(02.4375,QstateIM(3)) then
				char3IM <= "+02.4375";
			elsif QstateIM(3) = to_sfixed(02.5000,QstateIM(3)) then
				char3IM <= "+02.5000";
			elsif QstateIM(3) = to_sfixed(02.5625,QstateIM(3)) then
				char3IM <= "+02.5625";
			elsif QstateIM(3) = to_sfixed(02.6250,QstateIM(3)) then
				char3IM <= "+02.6250";
			elsif QstateIM(3) = to_sfixed(02.6875,QstateIM(3)) then
				char3IM <= "+02.6875";
			elsif QstateIM(3) = to_sfixed(02.7500,QstateIM(3)) then
				char3IM <= "+02.7500";
			elsif QstateIM(3) = to_sfixed(02.8125,QstateIM(3)) then
				char3IM <= "+02.8125";
			elsif QstateIM(3) = to_sfixed(02.8750,QstateIM(3)) then
				char3IM <= "+02.8750";
			elsif QstateIM(3) = to_sfixed(02.9375,QstateIM(3)) then
				char3IM <= "+02.9375";
			elsif QstateIM(3) = to_sfixed(03.0000,QstateIM(3)) then
				char3IM <= "+03.0000";
			elsif QstateIM(3) = to_sfixed(03.0625,QstateIM(3)) then
				char3IM <= "+03.0625";
			elsif QstateIM(3) = to_sfixed(03.1250,QstateIM(3)) then
				char3IM <= "+03.1250";
			elsif QstateIM(3) = to_sfixed(03.1875,QstateIM(3)) then
				char3IM <= "+03.1875";
			elsif QstateIM(3) = to_sfixed(03.2500,QstateIM(3)) then
				char3IM <= "+03.2500";
			elsif QstateIM(3) = to_sfixed(03.3125,QstateIM(3)) then
				char3IM <= "+03.3125";
			elsif QstateIM(3) = to_sfixed(03.3750,QstateIM(3)) then
				char3IM <= "+03.3750";
			elsif QstateIM(3) = to_sfixed(03.4375,QstateIM(3)) then
				char3IM <= "+03.4375";
			elsif QstateIM(3) = to_sfixed(03.5000,QstateIM(3)) then
				char3IM <= "+03.5000";
			elsif QstateIM(3) = to_sfixed(03.5625,QstateIM(3)) then
				char3IM <= "+03.5625";
			elsif QstateIM(3) = to_sfixed(03.6250,QstateIM(3)) then
				char3IM <= "+03.6250";
			elsif QstateIM(3) = to_sfixed(03.6875,QstateIM(3)) then
				char3IM <= "+03.6875";
			elsif QstateIM(3) = to_sfixed(03.7500,QstateIM(3)) then
				char3IM <= "+03.7500";
			elsif QstateIM(3) = to_sfixed(03.8125,QstateIM(3)) then
				char3IM <= "+03.8125";
			elsif QstateIM(3) = to_sfixed(03.8750,QstateIM(3)) then
				char3IM <= "+03.8750";
			elsif QstateIM(3) = to_sfixed(03.9375,QstateIM(3)) then
				char3IM <= "+03.9375";
			elsif QstateIM(3) = to_sfixed(04.0000,QstateIM(3)) then
				char3IM <= "+04.0000";
			elsif QstateIM(3) = to_sfixed(04.0625,QstateIM(3)) then
				char3IM <= "+04.0625";
			elsif QstateIM(3) = to_sfixed(04.1250,QstateIM(3)) then
				char3IM <= "+04.1250";
			elsif QstateIM(3) = to_sfixed(04.1875,QstateIM(3)) then
				char3IM <= "+04.1875";
			elsif QstateIM(3) = to_sfixed(04.2500,QstateIM(3)) then
				char3IM <= "+04.2500";
			elsif QstateIM(3) = to_sfixed(04.3125,QstateIM(3)) then
				char3IM <= "+04.3125";
			elsif QstateIM(3) = to_sfixed(04.3750,QstateIM(3)) then
				char3IM <= "+04.3750";
			elsif QstateIM(3) = to_sfixed(04.4375,QstateIM(3)) then
				char3IM <= "+04.4375";
			elsif QstateIM(3) = to_sfixed(04.5000,QstateIM(3)) then
				char3IM <= "+04.5000";
			elsif QstateIM(3) = to_sfixed(04.5625,QstateIM(3)) then
				char3IM <= "+04.5625";
			elsif QstateIM(3) = to_sfixed(04.6250,QstateIM(3)) then
				char3IM <= "+04.6250";
			elsif QstateIM(3) = to_sfixed(04.6875,QstateIM(3)) then
				char3IM <= "+04.6875";
			elsif QstateIM(3) = to_sfixed(04.7500,QstateIM(3)) then
				char3IM <= "+04.7500";
			elsif QstateIM(3) = to_sfixed(04.8125,QstateIM(3)) then
				char3IM <= "+04.8125";
			elsif QstateIM(3) = to_sfixed(04.8750,QstateIM(3)) then
				char3IM <= "+04.8750";
			elsif QstateIM(3) = to_sfixed(04.9375,QstateIM(3)) then
				char3IM <= "+04.9375";
			elsif QstateIM(3) = to_sfixed(05.0000,QstateIM(3)) then
				char3IM <= "+05.0000";
			elsif QstateIM(3) = to_sfixed(05.0625,QstateIM(3)) then
				char3IM <= "+05.0625";
			elsif QstateIM(3) = to_sfixed(05.1250,QstateIM(3)) then
				char3IM <= "+05.1250";
			elsif QstateIM(3) = to_sfixed(05.1875,QstateIM(3)) then
				char3IM <= "+05.1875";
			elsif QstateIM(3) = to_sfixed(05.2500,QstateIM(3)) then
				char3IM <= "+05.2500";
			elsif QstateIM(3) = to_sfixed(05.3125,QstateIM(3)) then
				char3IM <= "+05.3125";
			elsif QstateIM(3) = to_sfixed(05.3750,QstateIM(3)) then
				char3IM <= "+05.3750";
			elsif QstateIM(3) = to_sfixed(05.4375,QstateIM(3)) then
				char3IM <= "+05.4375";
			elsif QstateIM(3) = to_sfixed(05.5000,QstateIM(3)) then
				char3IM <= "+05.5000";
			elsif QstateIM(3) = to_sfixed(05.5625,QstateIM(3)) then
				char3IM <= "+05.5625";
			elsif QstateIM(3) = to_sfixed(05.6250,QstateIM(3)) then
				char3IM <= "+05.6250";
			elsif QstateIM(3) = to_sfixed(05.6875,QstateIM(3)) then
				char3IM <= "+05.6875";
			elsif QstateIM(3) = to_sfixed(05.7500,QstateIM(3)) then
				char3IM <= "+05.7500";
			elsif QstateIM(3) = to_sfixed(05.8125,QstateIM(3)) then
				char3IM <= "+05.8125";
			elsif QstateIM(3) = to_sfixed(05.8750,QstateIM(3)) then
				char3IM <= "+05.8750";
			elsif QstateIM(3) = to_sfixed(05.9375,QstateIM(3)) then
				char3IM <= "+05.9375";
			elsif QstateIM(3) = to_sfixed(06.0000,QstateIM(3)) then
				char3IM <= "+06.0000";
			elsif QstateIM(3) = to_sfixed(06.0625,QstateIM(3)) then
				char3IM <= "+06.0625";
			elsif QstateIM(3) = to_sfixed(06.1250,QstateIM(3)) then
				char3IM <= "+06.1250";
			elsif QstateIM(3) = to_sfixed(06.1875,QstateIM(3)) then
				char3IM <= "+06.1875";
			elsif QstateIM(3) = to_sfixed(06.2500,QstateIM(3)) then
				char3IM <= "+06.2500";
			elsif QstateIM(3) = to_sfixed(06.3125,QstateIM(3)) then
				char3IM <= "+06.3125";
			elsif QstateIM(3) = to_sfixed(06.3750,QstateIM(3)) then
				char3IM <= "+06.3750";
			elsif QstateIM(3) = to_sfixed(06.4375,QstateIM(3)) then
				char3IM <= "+06.4375";
			elsif QstateIM(3) = to_sfixed(06.5000,QstateIM(3)) then
				char3IM <= "+06.5000";
			elsif QstateIM(3) = to_sfixed(06.5625,QstateIM(3)) then
				char3IM <= "+06.5625";
			elsif QstateIM(3) = to_sfixed(06.6250,QstateIM(3)) then
				char3IM <= "+06.6250";
			elsif QstateIM(3) = to_sfixed(06.6875,QstateIM(3)) then
				char3IM <= "+06.6875";
			elsif QstateIM(3) = to_sfixed(06.7500,QstateIM(3)) then
				char3IM <= "+06.7500";
			elsif QstateIM(3) = to_sfixed(06.8125,QstateIM(3)) then
				char3IM <= "+06.8125";
			elsif QstateIM(3) = to_sfixed(06.8750,QstateIM(3)) then
				char3IM <= "+06.8750";
			elsif QstateIM(3) = to_sfixed(06.9375,QstateIM(3)) then
				char3IM <= "+06.9375";
			elsif QstateIM(3) = to_sfixed(07.0000,QstateIM(3)) then
				char3IM <= "+07.0000";
			elsif QstateIM(3) = to_sfixed(07.0625,QstateIM(3)) then
				char3IM <= "+07.0625";
			elsif QstateIM(3) = to_sfixed(07.1250,QstateIM(3)) then
				char3IM <= "+07.1250";
			elsif QstateIM(3) = to_sfixed(07.1875,QstateIM(3)) then
				char3IM <= "+07.1875";
			elsif QstateIM(3) = to_sfixed(07.2500,QstateIM(3)) then
				char3IM <= "+07.2500";
			elsif QstateIM(3) = to_sfixed(07.3125,QstateIM(3)) then
				char3IM <= "+07.3125";
			elsif QstateIM(3) = to_sfixed(07.3750,QstateIM(3)) then
				char3IM <= "+07.3750";
			elsif QstateIM(3) = to_sfixed(07.4375,QstateIM(3)) then
				char3IM <= "+07.4375";
			elsif QstateIM(3) = to_sfixed(07.5000,QstateIM(3)) then
				char3IM <= "+07.5000";
			elsif QstateIM(3) = to_sfixed(07.5625,QstateIM(3)) then
				char3IM <= "+07.5625";
			elsif QstateIM(3) = to_sfixed(07.6250,QstateIM(3)) then
				char3IM <= "+07.6250";
			elsif QstateIM(3) = to_sfixed(07.6875,QstateIM(3)) then
				char3IM <= "+07.6875";
			elsif QstateIM(3) = to_sfixed(07.7500,QstateIM(3)) then
				char3IM <= "+07.7500";
			elsif QstateIM(3) = to_sfixed(07.8125,QstateIM(3)) then
				char3IM <= "+07.8125";
			elsif QstateIM(3) = to_sfixed(07.8750,QstateIM(3)) then
				char3IM <= "+07.8750";
			elsif QstateIM(3) = to_sfixed(07.9375,QstateIM(3)) then
				char3IM <= "+07.9375";
			elsif QstateIM(3) = to_sfixed(08.0000,QstateIM(3)) then
				char3IM <= "+08.0000";
			elsif QstateIM(3) = to_sfixed(08.0625,QstateIM(3)) then
				char3IM <= "+08.0625";
			elsif QstateIM(3) = to_sfixed(08.1250,QstateIM(3)) then
				char3IM <= "+08.1250";
			elsif QstateIM(3) = to_sfixed(08.1875,QstateIM(3)) then
				char3IM <= "+08.1875";
			elsif QstateIM(3) = to_sfixed(08.2500,QstateIM(3)) then
				char3IM <= "+08.2500";
			elsif QstateIM(3) = to_sfixed(08.3125,QstateIM(3)) then
				char3IM <= "+08.3125";
			elsif QstateIM(3) = to_sfixed(08.3750,QstateIM(3)) then
				char3IM <= "+08.3750";
			elsif QstateIM(3) = to_sfixed(08.4375,QstateIM(3)) then
				char3IM <= "+08.4375";
			elsif QstateIM(3) = to_sfixed(08.5000,QstateIM(3)) then
				char3IM <= "+08.5000";
			elsif QstateIM(3) = to_sfixed(08.5625,QstateIM(3)) then
				char3IM <= "+08.5625";
			elsif QstateIM(3) = to_sfixed(08.6250,QstateIM(3)) then
				char3IM <= "+08.6250";
			elsif QstateIM(3) = to_sfixed(08.6875,QstateIM(3)) then
				char3IM <= "+08.6875";
			elsif QstateIM(3) = to_sfixed(08.7500,QstateIM(3)) then
				char3IM <= "+08.7500";
			elsif QstateIM(3) = to_sfixed(08.8125,QstateIM(3)) then
				char3IM <= "+08.8125";
			elsif QstateIM(3) = to_sfixed(08.8750,QstateIM(3)) then
				char3IM <= "+08.8750";
			elsif QstateIM(3) = to_sfixed(08.9375,QstateIM(3)) then
				char3IM <= "+08.9375";
			elsif QstateIM(3) = to_sfixed(09.0000,QstateIM(3)) then
				char3IM <= "+09.0000";
			elsif QstateIM(3) = to_sfixed(09.0625,QstateIM(3)) then
				char3IM <= "+09.0625";
			elsif QstateIM(3) = to_sfixed(09.1250,QstateIM(3)) then
				char3IM <= "+09.1250";
			elsif QstateIM(3) = to_sfixed(09.1875,QstateIM(3)) then
				char3IM <= "+09.1875";
			elsif QstateIM(3) = to_sfixed(09.2500,QstateIM(3)) then
				char3IM <= "+09.2500";
			elsif QstateIM(3) = to_sfixed(09.3125,QstateIM(3)) then
				char3IM <= "+09.3125";
			elsif QstateIM(3) = to_sfixed(09.3750,QstateIM(3)) then
				char3IM <= "+09.3750";
			elsif QstateIM(3) = to_sfixed(09.4375,QstateIM(3)) then
				char3IM <= "+09.4375";
			elsif QstateIM(3) = to_sfixed(09.5000,QstateIM(3)) then
				char3IM <= "+09.5000";
			elsif QstateIM(3) = to_sfixed(09.5625,QstateIM(3)) then
				char3IM <= "+09.5625";
			elsif QstateIM(3) = to_sfixed(09.6250,QstateIM(3)) then
				char3IM <= "+09.6250";
			elsif QstateIM(3) = to_sfixed(09.6875,QstateIM(3)) then
				char3IM <= "+09.6875";
			elsif QstateIM(3) = to_sfixed(09.7500,QstateIM(3)) then
				char3IM <= "+09.7500";
			elsif QstateIM(3) = to_sfixed(09.8125,QstateIM(3)) then
				char3IM <= "+09.8125";
			elsif QstateIM(3) = to_sfixed(09.8750,QstateIM(3)) then
				char3IM <= "+09.8750";
			elsif QstateIM(3) = to_sfixed(09.9375,QstateIM(3)) then
				char3IM <= "+09.9375";
			elsif QstateIM(3) = to_sfixed(10.0000,QstateIM(3)) then
				char3IM <= "+10.0000";
			elsif QstateIM(3) = to_sfixed(10.0625,QstateIM(3)) then
				char3IM <= "+10.0625";
			elsif QstateIM(3) = to_sfixed(10.1250,QstateIM(3)) then
				char3IM <= "+10.1250";
			elsif QstateIM(3) = to_sfixed(10.1875,QstateIM(3)) then
				char3IM <= "+10.1875";
			elsif QstateIM(3) = to_sfixed(10.2500,QstateIM(3)) then
				char3IM <= "+10.2500";
			elsif QstateIM(3) = to_sfixed(10.3125,QstateIM(3)) then
				char3IM <= "+10.3125";
			elsif QstateIM(3) = to_sfixed(10.3750,QstateIM(3)) then
				char3IM <= "+10.3750";
			elsif QstateIM(3) = to_sfixed(10.4375,QstateIM(3)) then
				char3IM <= "+10.4375";
			elsif QstateIM(3) = to_sfixed(10.5000,QstateIM(3)) then
				char3IM <= "+10.5000";
			elsif QstateIM(3) = to_sfixed(10.5625,QstateIM(3)) then
				char3IM <= "+10.5625";
			elsif QstateIM(3) = to_sfixed(10.6250,QstateIM(3)) then
				char3IM <= "+10.6250";
			elsif QstateIM(3) = to_sfixed(10.6875,QstateIM(3)) then
				char3IM <= "+10.6875";
			elsif QstateIM(3) = to_sfixed(10.7500,QstateIM(3)) then
				char3IM <= "+10.7500";
			elsif QstateIM(3) = to_sfixed(10.8125,QstateIM(3)) then
				char3IM <= "+10.8125";
			elsif QstateIM(3) = to_sfixed(10.8750,QstateIM(3)) then
				char3IM <= "+10.8750";
			elsif QstateIM(3) = to_sfixed(10.9375,QstateIM(3)) then
				char3IM <= "+10.9375";
			elsif QstateIM(3) = to_sfixed(11.0000,QstateIM(3)) then
				char3IM <= "+11.0000";
			elsif QstateIM(3) = to_sfixed(11.0625,QstateIM(3)) then
				char3IM <= "+11.0625";
			elsif QstateIM(3) = to_sfixed(11.1250,QstateIM(3)) then
				char3IM <= "+11.1250";
			elsif QstateIM(3) = to_sfixed(11.1875,QstateIM(3)) then
				char3IM <= "+11.1875";
			elsif QstateIM(3) = to_sfixed(11.2500,QstateIM(3)) then
				char3IM <= "+11.2500";
			elsif QstateIM(3) = to_sfixed(11.3125,QstateIM(3)) then
				char3IM <= "+11.3125";
			elsif QstateIM(3) = to_sfixed(11.3750,QstateIM(3)) then
				char3IM <= "+11.3750";
			elsif QstateIM(3) = to_sfixed(11.4375,QstateIM(3)) then
				char3IM <= "+11.4375";
			elsif QstateIM(3) = to_sfixed(11.5000,QstateIM(3)) then
				char3IM <= "+11.5000";
			elsif QstateIM(3) = to_sfixed(11.5625,QstateIM(3)) then
				char3IM <= "+11.5625";
			elsif QstateIM(3) = to_sfixed(11.6250,QstateIM(3)) then
				char3IM <= "+11.6250";
			elsif QstateIM(3) = to_sfixed(11.6875,QstateIM(3)) then
				char3IM <= "+11.6875";
			elsif QstateIM(3) = to_sfixed(11.7500,QstateIM(3)) then
				char3IM <= "+11.7500";
			elsif QstateIM(3) = to_sfixed(11.8125,QstateIM(3)) then
				char3IM <= "+11.8125";
			elsif QstateIM(3) = to_sfixed(11.8750,QstateIM(3)) then
				char3IM <= "+11.8750";
			elsif QstateIM(3) = to_sfixed(11.9375,QstateIM(3)) then
				char3IM <= "+11.9375";
			elsif QstateIM(3) = to_sfixed(12.0000,QstateIM(3)) then
				char3IM <= "+12.0000";
			elsif QstateIM(3) = to_sfixed(12.0625,QstateIM(3)) then
				char3IM <= "+12.0625";
			elsif QstateIM(3) = to_sfixed(12.1250,QstateIM(3)) then
				char3IM <= "+12.1250";
			elsif QstateIM(3) = to_sfixed(12.1875,QstateIM(3)) then
				char3IM <= "+12.1875";
			elsif QstateIM(3) = to_sfixed(12.2500,QstateIM(3)) then
				char3IM <= "+12.2500";
			elsif QstateIM(3) = to_sfixed(12.3125,QstateIM(3)) then
				char3IM <= "+12.3125";
			elsif QstateIM(3) = to_sfixed(12.3750,QstateIM(3)) then
				char3IM <= "+12.3750";
			elsif QstateIM(3) = to_sfixed(12.4375,QstateIM(3)) then
				char3IM <= "+12.4375";
			elsif QstateIM(3) = to_sfixed(12.5000,QstateIM(3)) then
				char3IM <= "+12.5000";
			elsif QstateIM(3) = to_sfixed(12.5625,QstateIM(3)) then
				char3IM <= "+12.5625";
			elsif QstateIM(3) = to_sfixed(12.6250,QstateIM(3)) then
				char3IM <= "+12.6250";
			elsif QstateIM(3) = to_sfixed(12.6875,QstateIM(3)) then
				char3IM <= "+12.6875";
			elsif QstateIM(3) = to_sfixed(12.7500,QstateIM(3)) then
				char3IM <= "+12.7500";
			elsif QstateIM(3) = to_sfixed(12.8125,QstateIM(3)) then
				char3IM <= "+12.8125";
			elsif QstateIM(3) = to_sfixed(12.8750,QstateIM(3)) then
				char3IM <= "+12.8750";
			elsif QstateIM(3) = to_sfixed(12.9375,QstateIM(3)) then
				char3IM <= "+12.9375";
			elsif QstateIM(3) = to_sfixed(13.0000,QstateIM(3)) then
				char3IM <= "+13.0000";
			elsif QstateIM(3) = to_sfixed(13.0625,QstateIM(3)) then
				char3IM <= "+13.0625";
			elsif QstateIM(3) = to_sfixed(13.1250,QstateIM(3)) then
				char3IM <= "+13.1250";
			elsif QstateIM(3) = to_sfixed(13.1875,QstateIM(3)) then
				char3IM <= "+13.1875";
			elsif QstateIM(3) = to_sfixed(13.2500,QstateIM(3)) then
				char3IM <= "+13.2500";
			elsif QstateIM(3) = to_sfixed(13.3125,QstateIM(3)) then
				char3IM <= "+13.3125";
			elsif QstateIM(3) = to_sfixed(13.3750,QstateIM(3)) then
				char3IM <= "+13.3750";
			elsif QstateIM(3) = to_sfixed(13.4375,QstateIM(3)) then
				char3IM <= "+13.4375";
			elsif QstateIM(3) = to_sfixed(13.5000,QstateIM(3)) then
				char3IM <= "+13.5000";
			elsif QstateIM(3) = to_sfixed(13.5625,QstateIM(3)) then
				char3IM <= "+13.5625";
			elsif QstateIM(3) = to_sfixed(13.6250,QstateIM(3)) then
				char3IM <= "+13.6250";
			elsif QstateIM(3) = to_sfixed(13.6875,QstateIM(3)) then
				char3IM <= "+13.6875";
			elsif QstateIM(3) = to_sfixed(13.7500,QstateIM(3)) then
				char3IM <= "+13.7500";
			elsif QstateIM(3) = to_sfixed(13.8125,QstateIM(3)) then
				char3IM <= "+13.8125";
			elsif QstateIM(3) = to_sfixed(13.8750,QstateIM(3)) then
				char3IM <= "+13.8750";
			elsif QstateIM(3) = to_sfixed(13.9375,QstateIM(3)) then
				char3IM <= "+13.9375";
			elsif QstateIM(3) = to_sfixed(14.0000,QstateIM(3)) then
				char3IM <= "+14.0000";
			elsif QstateIM(3) = to_sfixed(14.0625,QstateIM(3)) then
				char3IM <= "+14.0625";
			elsif QstateIM(3) = to_sfixed(14.1250,QstateIM(3)) then
				char3IM <= "+14.1250";
			elsif QstateIM(3) = to_sfixed(14.1875,QstateIM(3)) then
				char3IM <= "+14.1875";
			elsif QstateIM(3) = to_sfixed(14.2500,QstateIM(3)) then
				char3IM <= "+14.2500";
			elsif QstateIM(3) = to_sfixed(14.3125,QstateIM(3)) then
				char3IM <= "+14.3125";
			elsif QstateIM(3) = to_sfixed(14.3750,QstateIM(3)) then
				char3IM <= "+14.3750";
			elsif QstateIM(3) = to_sfixed(14.4375,QstateIM(3)) then
				char3IM <= "+14.4375";
			elsif QstateIM(3) = to_sfixed(14.5000,QstateIM(3)) then
				char3IM <= "+14.5000";
			elsif QstateIM(3) = to_sfixed(14.5625,QstateIM(3)) then
				char3IM <= "+14.5625";
			elsif QstateIM(3) = to_sfixed(14.6250,QstateIM(3)) then
				char3IM <= "+14.6250";
			elsif QstateIM(3) = to_sfixed(14.6875,QstateIM(3)) then
				char3IM <= "+14.6875";
			elsif QstateIM(3) = to_sfixed(14.7500,QstateIM(3)) then
				char3IM <= "+14.7500";
			elsif QstateIM(3) = to_sfixed(14.8125,QstateIM(3)) then
				char3IM <= "+14.8125";
			elsif QstateIM(3) = to_sfixed(14.8750,QstateIM(3)) then
				char3IM <= "+14.8750";
			elsif QstateIM(3) = to_sfixed(14.9375,QstateIM(3)) then
				char3IM <= "+14.9375";
			elsif QstateIM(3) = to_sfixed(15.0000,QstateIM(3)) then
				char3IM <= "+15.0000";
			elsif QstateIM(3) = to_sfixed(15.0625,QstateIM(3)) then
				char3IM <= "+15.0625";
			elsif QstateIM(3) = to_sfixed(15.1250,QstateIM(3)) then
				char3IM <= "+15.1250";
			elsif QstateIM(3) = to_sfixed(15.1875,QstateIM(3)) then
				char3IM <= "+15.1875";
			elsif QstateIM(3) = to_sfixed(15.2500,QstateIM(3)) then
				char3IM <= "+15.2500";
			elsif QstateIM(3) = to_sfixed(15.3125,QstateIM(3)) then
				char3IM <= "+15.3125";
			elsif QstateIM(3) = to_sfixed(15.3750,QstateIM(3)) then
				char3IM <= "+15.3750";
			elsif QstateIM(3) = to_sfixed(15.4375,QstateIM(3)) then
				char3IM <= "+15.4375";
			elsif QstateIM(3) = to_sfixed(15.5000,QstateIM(3)) then
				char3IM <= "+15.5000";
			elsif QstateIM(3) = to_sfixed(15.5625,QstateIM(3)) then
				char3IM <= "+15.5625";
			elsif QstateIM(3) = to_sfixed(15.6250,QstateIM(3)) then
				char3IM <= "+15.6250";
			elsif QstateIM(3) = to_sfixed(15.6875,QstateIM(3)) then
				char3IM <= "+15.6875";
			elsif QstateIM(3) = to_sfixed(15.7500,QstateIM(3)) then
				char3IM <= "+15.7500";
			elsif QstateIM(3) = to_sfixed(15.8125,QstateIM(3)) then
				char3IM <= "+15.8125";
			elsif QstateIM(3) = to_sfixed(15.8750,QstateIM(3)) then
				char3IM <= "+15.8750";
			elsif QstateIM(3) = to_sfixed(15.9375,QstateIM(3)) then
				char3IM <= "+15.9375";
			end if;
		state_next <= Stitch;
		
		when Stitch =>
			Output(1 to 8) <= char0RE; --& char0IM & char1RE & char1IM & char2RE & char2IM & char3RE & char3IM ;
			Output(9 to 16) <= char0IM;
			Output(17 to 24) <= char1RE;
			Output(25 to 32) <= char1IM;
			Output(33 to 40) <= char2RE;
			Output(41 to 48) <= char2IM;
			Output(49 to 56) <= char3RE;
			Output(57 to 64) <= char3IM;
			state_next <= finish;				
			
		when finish =>
			finished <= '1';

		end case;
		end process QFT;
end compute;