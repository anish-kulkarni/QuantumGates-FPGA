library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.MATH_REAL.ALL;


library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
use ieee_proposed.float_pkg.all;


------------------------
-- ENTITY DECLARATION --
------------------------

entity float_mult is
	port(
			--in1 : in sfixed(1 downto -2);
			--in2 : in sfixed(1 downto -2);
			clk : in std_logic;
			product : out ufixed(3 downto -4);
			inter_state : in std_logic:= '0'
	);
end entity;

-------------------------
-- ARCHITECTURE DECLARATION --
-------------------------

architecture behave of float_mult is
signal temp : ufixed(3 downto -4);
--signal temp2 : ufixed(3 downto -4);
signal in1 : ufixed(1 downto -2):="1001"; --in1 = 2.25
signal in2 : ufixed(1 downto -2):="1101"; --in2 = 3.25
--signal result :string(1 to 9);
begin
process(clk)
	begin
	
		temp <= in1*in2; -- product = 8.75 (in decimal) = 1000.1100
		

			product <= temp;
		
		
	end process;	
	
	
--		conv : process(temp, inter_state) 
--		begin
--			
--				if temp = "00000000" then
--					result <= "00.0000";
--				elsif temp = "00000001" then
--					result <= "00.0625";
--				elsif temp = "00000010" then
--					result <= "00.1250";
--				elsif temp = "00000011" then
--					result <= "00.1875";
--				elsif temp = "00000100" then
--					result <= "00.2500";
--				elsif temp = "00000101" then
--					result <= "00.3125";
--				elsif temp = "00000110" then
--					result <= "00.3750";
--				elsif temp = "00000111" then
--					result <= "00.4375";
--				elsif temp = "00001000" then
--					result <= "00.5000";
--				elsif temp = "00001001" then
--					result <= "00.5625";
--				elsif temp = "00001010" then
--					result <= "00.6250";
--				elsif temp = "00001011" then
--					result <= "00.6875";
--				elsif temp = "00001100" then
--					result <= "00.7500";
--				elsif temp = "00001101" then
--					result <= "00.8125";
--				elsif temp = "00001110" then
--					result <= "00.8750";
--				elsif temp = "00001111" then
--					result <= "00.9375";
--				elsif temp = "00010000" then
--					result <= "01.0000";
--				elsif temp = "00010001" then
--					result <= "01.0625";
--				elsif temp = "00010010" then
--					result <= "01.1250";
--				elsif temp = "00010011" then
--					result <= "01.1875";
--				elsif temp = "00010100" then
--					result <= "01.2500";
--				elsif temp = "00010101" then
--					result <= "01.3125";
--				elsif temp = "00010110" then
--					result <= "01.3750";
--				elsif temp = "00010111" then
--					result <= "01.4375";
--				elsif temp = "00011000" then
--					result <= "01.5000";
--				elsif temp = "00011001" then
--					result <= "01.5625";
--				elsif temp = "00011010" then
--					result <= "01.6250";
--				elsif temp = "00011011" then
--					result <= "01.6875";
--				elsif temp = "00011100" then
--					result <= "01.7500";
--				elsif temp = "00011101" then
--					result <= "01.8125";
--				elsif temp = "00011110" then
--					result <= "01.8750";
--				elsif temp = "00011111" then
--					result <= "01.9375";
--				elsif temp = "00100000" then
--					result <= "02.0000";
--				elsif temp = "00100001" then
--					result <= "02.0625";
--				elsif temp = "00100010" then
--					result <= "02.1250";
--				elsif temp = "00100011" then
--					result <= "02.1875";
--				elsif temp = "00100100" then
--					result <= "02.2500";
--				elsif temp = "00100101" then
--					result <= "02.3125";
--				elsif temp = "00100110" then
--					result <= "02.3750";
--				elsif temp = "00100111" then
--					result <= "02.4375";
--				elsif temp = "00101000" then
--					result <= "02.5000";
--				elsif temp = "00101001" then
--					result <= "02.5625";
--				elsif temp = "00101010" then
--					result <= "02.6250";
--				elsif temp = "00101011" then
--					result <= "02.6875";
--				elsif temp = "00101100" then
--					result <= "02.7500";
--				elsif temp = "00101101" then
--					result <= "02.8125";
--				elsif temp = "00101110" then
--					result <= "02.8750";
--				elsif temp = "00101111" then
--					result <= "02.9375";
--				elsif temp = "00110000" then
--					result <= "03.0000";
--				elsif temp = "00110001" then
--					result <= "03.0625";
--				elsif temp = "00110010" then
--					result <= "03.1250";
--				elsif temp = "00110011" then
--					result <= "03.1875";
--				elsif temp = "00110100" then
--					result <= "03.2500";
--				elsif temp = "00110101" then
--					result <= "03.3125";
--				elsif temp = "00110110" then
--					result <= "03.3750";
--				elsif temp = "00110111" then
--					result <= "03.4375";
--				elsif temp = "00111000" then
--					result <= "03.5000";
--				elsif temp = "00111001" then
--					result <= "03.5625";
--				elsif temp = "00111010" then
--					result <= "03.6250";
--				elsif temp = "00111011" then
--					result <= "03.6875";
--				elsif temp = "00111100" then
--					result <= "03.7500";
--				elsif temp = "00111101" then
--					result <= "03.8125";
--				elsif temp = "00111110" then
--					result <= "03.8750";
--				elsif temp = "00111111" then
--					result <= "03.9375";
--				elsif temp = "01000000" then
--					result <= "04.0000";
--				elsif temp = "01000001" then
--					result <= "04.0625";
--				elsif temp = "01000010" then
--					result <= "04.1250";
--				elsif temp = "01000011" then
--					result <= "04.1875";
--				elsif temp = "01000100" then
--					result <= "04.2500";
--				elsif temp = "01000101" then
--					result <= "04.3125";
--				elsif temp = "01000110" then
--					result <= "04.3750";
--				elsif temp = "01000111" then
--					result <= "04.4375";
--				elsif temp = "01001000" then
--					result <= "04.5000";
--				elsif temp = "01001001" then
--					result <= "04.5625";
--				elsif temp = "01001010" then
--					result <= "04.6250";
--				elsif temp = "01001011" then
--					result <= "04.6875";
--				elsif temp = "01001100" then
--					result <= "04.7500";
--				elsif temp = "01001101" then
--					result <= "04.8125";
--				elsif temp = "01001110" then
--					result <= "04.8750";
--				elsif temp = "01001111" then
--					result <= "04.9375";
--				elsif temp = "01010000" then
--					result <= "05.0000";
--				elsif temp = "01010001" then
--					result <= "05.0625";
--				elsif temp = "01010010" then
--					result <= "05.1250";
--				elsif temp = "01010011" then
--					result <= "05.1875";
--				elsif temp = "01010100" then
--					result <= "05.2500";
--				elsif temp = "01010101" then
--					result <= "05.3125";
--				elsif temp = "01010110" then
--					result <= "05.3750";
--				elsif temp = "01010111" then
--					result <= "05.4375";
--				elsif temp = "01011000" then
--					result <= "05.5000";
--				elsif temp = "01011001" then
--					result <= "05.5625";
--				elsif temp = "01011010" then
--					result <= "05.6250";
--				elsif temp = "01011011" then
--					result <= "05.6875";
--				elsif temp = "01011100" then
--					result <= "05.7500";
--				elsif temp = "01011101" then
--					result <= "05.8125";
--				elsif temp = "01011110" then
--					result <= "05.8750";
--				elsif temp = "01011111" then
--					result <= "05.9375";
--				elsif temp = "01100000" then
--					result <= "06.0000";
--				elsif temp = "01100001" then
--					result <= "06.0625";
--				elsif temp = "01100010" then
--					result <= "06.1250";
--				elsif temp = "01100011" then
--					result <= "06.1875";
--				elsif temp = "01100100" then
--					result <= "06.2500";
--				elsif temp = "01100101" then
--					result <= "06.3125";
--				elsif temp = "01100110" then
--					result <= "06.3750";
--				elsif temp = "01100111" then
--					result <= "06.4375";
--				elsif temp = "01101000" then
--					result <= "06.5000";
--				elsif temp = "01101001" then
--					result <= "06.5625";
--				elsif temp = "01101010" then
--					result <= "06.6250";
--				elsif temp = "01101011" then
--					result <= "06.6875";
--				elsif temp = "01101100" then
--					result <= "06.7500";
--				elsif temp = "01101101" then
--					result <= "06.8125";
--				elsif temp = "01101110" then
--					result <= "06.8750";
--				elsif temp = "01101111" then
--					result <= "06.9375";
--				elsif temp = "01110000" then
--					result <= "07.0000";
--				elsif temp = "01110001" then
--					result <= "07.0625";
--				elsif temp = "01110010" then
--					result <= "07.1250";
--				elsif temp = "01110011" then
--					result <= "07.1875";
--				elsif temp = "01110100" then
--					result <= "07.2500";
--				elsif temp = "01110101" then
--					result <= "07.3125";
--				elsif temp = "01110110" then
--					result <= "07.3750";
--				elsif temp = "01110111" then
--					result <= "07.4375";
--				elsif temp = "01111000" then
--					result <= "07.5000";
--				elsif temp = "01111001" then
--					result <= "07.5625";
--				elsif temp = "01111010" then
--					result <= "07.6250";
--				elsif temp = "01111011" then
--					result <= "07.6875";
--				elsif temp = "01111100" then
--					result <= "07.7500";
--				elsif temp = "01111101" then
--					result <= "07.8125";
--				elsif temp = "01111110" then
--					result <= "07.8750";
--				elsif temp = "01111111" then
--					result <= "07.9375";
--				elsif temp = "10000000" then
--					result <= "08.0000";
--				elsif temp = "10000001" then
--					result <= "08.0625";
--				elsif temp = "10000010" then
--					result <= "08.1250";
--				elsif temp = "10000011" then
--					result <= "08.1875";
--				elsif temp = "10000100" then
--					result <= "08.2500";
--				elsif temp = "10000101" then
--					result <= "08.3125";
--				elsif temp = "10000110" then
--					result <= "08.3750";
--				elsif temp = "10000111" then
--					result <= "08.4375";
--				elsif temp = "10001000" then
--					result <= "08.5000";
--				elsif temp = "10001001" then
--					result <= "08.5625";
--				elsif temp = "10001010" then
--					result <= "08.6250";
--				elsif temp = "10001011" then
--					result <= "08.6875";
--				elsif temp = "10001100" then
--					result <= "08.7500";
--				elsif temp = "10001101" then
--					result <= "08.8125";
--				elsif temp = "10001110" then
--					result <= "08.8750";
--				elsif temp = "10001111" then
--					result <= "08.9375";
--				elsif temp = "10010000" then
--					result <= "09.0000";
--				elsif temp = "10010001" then
--					result <= "09.0625";
--				elsif temp = "10010010" then
--					result <= "09.1250";
--				elsif temp = "10010011" then
--					result <= "09.1875";
--				elsif temp = "10010100" then
--					result <= "09.2500";
--				elsif temp = "10010101" then
--					result <= "09.3125";
--				elsif temp = "10010110" then
--					result <= "09.3750";
--				elsif temp = "10010111" then
--					result <= "09.4375";
--				elsif temp = "10011000" then
--					result <= "09.5000";
--				elsif temp = "10011001" then
--					result <= "09.5625";
--				elsif temp = "10011010" then
--					result <= "09.6250";
--				elsif temp = "10011011" then
--					result <= "09.6875";
--				elsif temp = "10011100" then
--					result <= "09.7500";
--				elsif temp = "10011101" then
--					result <= "09.8125";
--				elsif temp = "10011110" then
--					result <= "09.8750";
--				elsif temp = "10011111" then
--					result <= "09.9375";
--				elsif temp = "10100000" then
--					result <= "10.0000";
--				elsif temp = "10100001" then
--					result <= "10.0625";
--				elsif temp = "10100010" then
--					result <= "10.1250";
--				elsif temp = "10100011" then
--					result <= "10.1875";
--				elsif temp = "10100100" then
--					result <= "10.2500";
--				elsif temp = "10100101" then
--					result <= "10.3125";
--				elsif temp = "10100110" then
--					result <= "10.3750";
--				elsif temp = "10100111" then
--					result <= "10.4375";
--				elsif temp = "10101000" then
--					result <= "10.5000";
--				elsif temp = "10101001" then
--					result <= "10.5625";
--				elsif temp = "10101010" then
--					result <= "10.6250";
--				elsif temp = "10101011" then
--					result <= "10.6875";
--				elsif temp = "10101100" then
--					result <= "10.7500";
--				elsif temp = "10101101" then
--					result <= "10.8125";
--				elsif temp = "10101110" then
--					result <= "10.8750";
--				elsif temp = "10101111" then
--					result <= "10.9375";
--				elsif temp = "10110000" then
--					result <= "11.0000";
--				elsif temp = "10110001" then
--					result <= "11.0625";
--				elsif temp = "10110010" then
--					result <= "11.1250";
--				elsif temp = "10110011" then
--					result <= "11.1875";
--				elsif temp = "10110100" then
--					result <= "11.2500";
--				elsif temp = "10110101" then
--					result <= "11.3125";
--				elsif temp = "10110110" then
--					result <= "11.3750";
--				elsif temp = "10110111" then
--					result <= "11.4375";
--				elsif temp = "10111000" then
--					result <= "11.5000";
--				elsif temp = "10111001" then
--					result <= "11.5625";
--				elsif temp = "10111010" then
--					result <= "11.6250";
--				elsif temp = "10111011" then
--					result <= "11.6875";
--				elsif temp = "10111100" then
--					result <= "11.7500";
--				elsif temp = "10111101" then
--					result <= "11.8125";
--				elsif temp = "10111110" then
--					result <= "11.8750";
--				elsif temp = "10111111" then
--					result <= "11.9375";
--				elsif temp = "11000000" then
--					result <= "12.0000";
--				elsif temp = "11000001" then
--					result <= "12.0625";
--				elsif temp = "11000010" then
--					result <= "12.1250";
--				elsif temp = "11000011" then
--					result <= "12.1875";
--				elsif temp = "11000100" then
--					result <= "12.2500";
--				elsif temp = "11000101" then
--					result <= "12.3125";
--				elsif temp = "11000110" then
--					result <= "12.3750";
--				elsif temp = "11000111" then
--					result <= "12.4375";
--				elsif temp = "11001000" then
--					result <= "12.5000";
--				elsif temp = "11001001" then
--					result <= "12.5625";
--				elsif temp = "11001010" then
--					result <= "12.6250";
--				elsif temp = "11001011" then
--					result <= "12.6875";
--				elsif temp = "11001100" then
--					result <= "12.7500";
--				elsif temp = "11001101" then
--					result <= "12.8125";
--				elsif temp = "11001110" then
--					result <= "12.8750";
--				elsif temp = "11001111" then
--					result <= "12.9375";
--				elsif temp = "11010000" then
--					result <= "13.0000";
--				elsif temp = "11010001" then
--					result <= "13.0625";
--				elsif temp = "11010010" then
--					result <= "13.1250";
--				elsif temp = "11010011" then
--					result <= "13.1875";
--				elsif temp = "11010100" then
--					result <= "13.2500";
--				elsif temp = "11010101" then
--					result <= "13.3125";
--				elsif temp = "11010110" then
--					result <= "13.3750";
--				elsif temp = "11010111" then
--					result <= "13.4375";
--				elsif temp = "11011000" then
--					result <= "13.5000";
--				elsif temp = "11011001" then
--					result <= "13.5625";
--				elsif temp = "11011010" then
--					result <= "13.6250";
--				elsif temp = "11011011" then
--					result <= "13.6875";
--				elsif temp = "11011100" then
--					result <= "13.7500";
--				elsif temp = "11011101" then
--					result <= "13.8125";
--				elsif temp = "11011110" then
--					result <= "13.8750";
--				elsif temp = "11011111" then
--					result <= "13.9375";
--				elsif temp = "11100000" then
--					result <= "14.0000";
--				elsif temp = "11100001" then
--					result <= "14.0625";
--				elsif temp = "11100010" then
--					result <= "14.1250";
--				elsif temp = "11100011" then
--					result <= "14.1875";
--				elsif temp = "11100100" then
--					result <= "14.2500";
--				elsif temp = "11100101" then
--					result <= "14.3125";
--				elsif temp = "11100110" then
--					result <= "14.3750";
--				elsif temp = "11100111" then
--					result <= "14.4375";
--				elsif temp = "11101000" then
--					result <= "14.5000";
--				elsif temp = "11101001" then
--					result <= "14.5625";
--				elsif temp = "11101010" then
--					result <= "14.6250";
--				elsif temp = "11101011" then
--					result <= "14.6875";
--				elsif temp = "11101100" then
--					result <= "14.7500";
--				elsif temp = "11101101" then
--					result <= "14.8125";
--				elsif temp = "11101110" then
--					result <= "14.8750";
--				elsif temp = "11101111" then
--					result <= "14.9375";
--				elsif temp = "11110000" then
--					result <= "15.0000";
--				elsif temp = "11110001" then
--					result <= "15.0625";
--				elsif temp = "11110010" then
--					result <= "15.1250";
--				elsif temp = "11110011" then
--					result <= "15.1875";
--				elsif temp = "11110100" then
--					result <= "15.2500";
--				elsif temp = "11110101" then
--					result <= "15.3125";
--				elsif temp = "11110110" then
--					result <= "15.3750";
--				elsif temp = "11110111" then
--					result <= "15.4375";
--				elsif temp = "11111000" then
--					result <= "15.5000";
--				elsif temp = "11111001" then
--					result <= "15.5625";
--				elsif temp = "11111010" then
--					result <= "15.6250";
--				elsif temp = "11111011" then
--					result <= "15.6875";
--				elsif temp = "11111100" then
--					result <= "15.7500";
--				elsif temp = "11111101" then
--					result <= "15.8125";
--				elsif temp = "11111110" then
--					result <= "15.8750";
--				elsif temp = "11111111" then
--					result <= "15.9375";
--				end if;
--
--		end process conv;
--			
			
		--end if;
	--end process;
	
end behave;